module macro_args_sub();
	`BAR(0)
endmodule
