module test;

reg [7:0] value, value;

endmodule
