module test();
// wire r;
a ua ( .r ( !r ));
endmodule

module a ( r );
input  r;
endmodule
