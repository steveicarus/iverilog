/*
 * Copyright (c) 1998-2000 Andrei Purdea (andrei@purdea.ro)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 */

// This test checks that returning from a void function works correctly.
module main;
  int res = 123;
  function void bla();
    int i;
    for (i=0;i<10;i=i+1) begin
        res = i;
        $display("loop %d", i);
        if (i == 5)
        begin
            return;
        end
    end
  endfunction
  initial begin
    bla();
    if (res == 5) begin
      $display("PASS");
    end else begin
      $display("FAIL");
    end
  end
endmodule
