module top;
  initial $display("The following should be a single percent: %");
endmodule
