`include "pr2215342_inc.v" // Include a file

module top;
  initial $display("PASSED");
endmodule
