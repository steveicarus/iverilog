module m;
  task t1;
    input make_me_crash i;
    begin
    end
  endtask
  task t2;
    input integer i;
    begin
    end
  endtask
endmodule
