module test;
    initial begin
	$display("Error: \"FloatTest.bsv\", line 234, column 24: (R0001)\n  Mutually exclusive rules (from the ME sets [RL_action_l234c24] and\n  [RL_action_l235c24, RL_action_l236c24, RL_action_l237c24, RL_action_l238c24,\n  RL_action_l239c24, RL_action_l240c24, RL_action_l241c24, RL_action_l242c24,\n  RL_action_l243c24, RL_action_l244c24, RL_action_l245c24, RL_action_l246c24,\n  RL_action_l247c24, RL_action_l248c24, RL_action_l249c24, RL_action_l250c24,\n  RL_action_l251c24, RL_action_l252c24, RL_action_l253c24, RL_action_l255c24,\n  RL_action_l256c24, RL_action_l257c24, RL_action_l258c24, RL_action_l259c24,\n  RL_action_l260c24, RL_action_l261c24, RL_action_l262c24, RL_action_l263c24,\n  RL_action_l264c24, RL_action_l265c24, RL_action_l266c24, RL_action_l267c24,\n  RL_action_l268c24, RL_action_l269c24, RL_action_l270c24, RL_action_l271c24,\n  RL_action_l272c24, RL_action_l273c24, RL_action_l274c24, RL_action_l276c24,\n  RL_action_l277c24, RL_action_l278c24, RL_action_l279c24, RL_action_l280c24,\n  RL_action_l281c24, RL_action_l282c24, RL_action_l283c24, RL_action_l284c24,\n  RL_action_l285c24, RL_action_l286c24, RL_action_l287c24, RL_action_l288c24,\n  RL_action_l289c24, RL_action_l290c24, RL_action_l291c24, RL_action_l292c24,\n  RL_action_l293c24, RL_action_l294c24, RL_action_l295c24, RL_action_l297c24,\n  RL_action_l298c24, RL_action_l299c24, RL_action_l300c24, RL_action_l301c24,\n  RL_action_l302c24, RL_action_l303c24, RL_action_l304c24, RL_action_l305c24,\n  RL_action_l306c24, RL_action_l307c24, RL_action_l308c24, RL_action_l309c24,\n  RL_action_l310c24, RL_action_l311c24, RL_action_l312c24, RL_action_l313c24,\n  RL_action_l314c24, RL_action_l315c24, RL_action_l316c24, RL_action_l318c24,\n  RL_action_l319c24, RL_action_l320c24, RL_action_l321c24, RL_action_l322c24,\n  RL_action_l323c24, RL_action_l324c24, RL_action_l326c24, RL_action_l327c24,\n  RL_action_l328c24, RL_action_l329c24, RL_action_l330c24, RL_action_l331c24,\n  RL_action_l332c24, RL_action_l333c24, RL_action_l334c24, RL_action_l335c24,\n  RL_action_l336c24, RL_action_l337c24, RL_action_l338c24, RL_action_l339c24,\n  RL_action_l340c24, RL_action_l341c24, RL_action_l342c24, RL_action_l343c24,\n  RL_action_l344c24, RL_action_l345c24, RL_action_l348c18, RL_action_l353c22,\n  RL_action_l354c22, RL_action_l355c22, RL_action_l356c22, RL_action_l357c22,\n  RL_action_l358c22, RL_action_l359c22, RL_action_l360c22, RL_action_l361c22,\n  RL_action_l362c22, RL_action_l363c22, RL_action_l364c22, RL_action_l365c22,\n  RL_action_l366c22, RL_action_l367c22, RL_action_l368c22, RL_action_l369c22,\n  RL_action_l370c22, RL_action_l371c22, RL_action_l372c22, RL_action_l374c22,\n  RL_action_l376c22, RL_action_l377c22, RL_action_l378c22, RL_action_l379c22,\n  RL_action_l381c22, RL_action_l383c22, RL_action_l384c22, RL_action_l386c22,\n  RL_action_l387c22, RL_action_l390c18, RL_action_l395c23, RL_action_l396c23,\n  RL_action_l398c23, RL_action_l399c23, RL_action_l400c23, RL_action_l401c23,\n  RL_action_l402c23, RL_action_l403c23, RL_action_l404c23, RL_action_l405c23,\n  RL_action_l406c23, RL_action_l407c23, RL_action_l408c23, RL_action_l409c23,\n  RL_action_l410c23, RL_action_l411c23, RL_action_l412c23, RL_action_l413c23,\n  RL_action_l414c23, RL_action_l415c23, RL_action_l416c23, RL_action_l417c23,\n  RL_action_l419c23, RL_action_l420c23, RL_action_l421c23, RL_action_l422c23,\n  RL_action_l423c23, RL_action_l424c23, RL_action_l425c23, RL_action_l426c23,\n  RL_action_l427c23, RL_action_l428c23, RL_action_l429c23, RL_action_l430c23,\n  RL_action_l431c23, RL_action_l432c23, RL_action_l433c23, RL_action_l434c23,\n  RL_action_l435c23, RL_action_l436c23, RL_action_l437c23, RL_action_l438c23,\n  RL_action_l441c18, RL_action_l446c28, RL_action_l447c28, RL_action_l448c28,\n  RL_action_l449c28, RL_action_l450c28, RL_action_l451c28, RL_action_l452c28,\n  RL_action_l453c28, RL_action_l455c28, RL_action_l456c28, RL_action_l457c28,\n  RL_action_l458c28, RL_action_l459c28, RL_action_l460c28, RL_action_l461c28,\n  RL_action_l462c28, RL_action_l463c28, RL_action_l464c28, RL_action_l465c28,\n  RL_action_l466c28, RL_action_l467c28, RL_action_l468c28, RL_action_l469c28,\n  RL_action_l470c28, RL_action_l471c28, RL_action_l472c28, RL_action_l473c28,\n  RL_action_l474c28, RL_action_l475c28, RL_action_l476c28, RL_action_l478c28,\n  RL_action_l479c28, RL_action_l481c28, RL_action_l484c18, RL_action_l489c21,\n  RL_action_l490c21, RL_action_l491c21, RL_action_l492c21, RL_action_l493c21,\n  RL_action_l494c21, RL_action_l495c21, RL_action_l496c21, RL_action_l497c21,\n  RL_action_l498c21, RL_action_l499c21, RL_action_l500c21, RL_action_l501c21,\n  RL_action_l502c21, RL_action_l503c21, RL_action_l504c21, RL_action_l505c21,\n  RL_action_l506c21, RL_action_l507c21, RL_action_l508c21, RL_action_l509c21,\n  RL_action_l510c21, RL_action_l512c21, RL_action_l513c21, RL_action_l514c21,\n  RL_action_l515c21, RL_action_l516c21, RL_action_l517c21, RL_action_l518c21,\n  RL_action_l519c21, RL_action_l520c21, RL_action_l521c21, RL_action_l522c21,\n  RL_action_l523c21, RL_action_l524c21, RL_action_l525c21, RL_action_l526c21,\n  RL_action_l527c21, RL_action_l528c21, RL_action_l529c21, RL_action_l530c21,\n  RL_action_l531c21, RL_action_l533c26, RL_action_l534c26, RL_action_l535c26,\n  RL_action_l536c26, RL_action_l537c26, RL_action_l538c26, RL_action_l539c26,\n  RL_action_l540c26, RL_action_l542c26, RL_action_l543c26, RL_action_l544c26,\n  RL_action_l545c26, RL_action_l546c26, RL_action_l547c26, RL_action_l548c26,\n  RL_action_l549c26, RL_action_l550c26, RL_action_l551c26, RL_action_l552c26,\n  RL_action_l553c26, RL_action_l554c26, RL_action_l555c26, RL_action_l556c26,\n  RL_action_l557c26, RL_action_l558c26, RL_action_l559c26, RL_action_l560c26,\n  RL_action_l561c26, RL_action_l562c26, RL_action_l563c26, RL_action_l565c26,\n  RL_action_l566c26, RL_action_l568c26, RL_action_l570c21, RL_action_l572c21,\n  RL_action_l574c26, RL_action_l576c26, RL_action_l577c26, RL_action_l579c26,\n  RL_action_l582c18, RL_action_l587c28, RL_action_l588c28, RL_action_l589c28,\n  RL_action_l590c28, RL_action_l591c28, RL_action_l592c28, RL_action_l593c28,\n  RL_action_l594c28, RL_action_l595c28, RL_action_l596c28, RL_action_l597c28,\n  RL_action_l598c28, RL_action_l599c28, RL_action_l600c28, RL_action_l601c28,\n  RL_action_l602c28, RL_action_l603c28, RL_action_l604c28, RL_action_l605c28,\n  RL_action_l606c28, RL_action_l607c28, RL_action_l609c28, RL_action_l610c28,\n  RL_action_l611c28, RL_action_l613c28, RL_action_l614c28, RL_action_l615c28,\n  RL_action_l616c28, RL_action_l617c28, RL_action_l618c28, RL_action_l619c28,\n  RL_action_l621c28, RL_action_l622c28, RL_action_l623c28, RL_action_l624c28,\n  RL_action_l625c28, RL_action_l626c28, RL_action_l627c28, RL_action_l628c28,\n  RL_action_l629c28, RL_action_l630c28, RL_action_l631c28, RL_action_l632c28,\n  RL_action_l633c28, RL_action_l634c28, RL_action_l635c28, RL_action_l636c28,\n  RL_action_l637c28, RL_action_l638c28, RL_action_l639c28, RL_action_l645c18,\n  RL_action_l647c7] ) fired in the same clock cycle.\nPASSED");
    end
endmodule
