/* )* */
/* (* /* *) */
module test();
initial $display("PASSED");
endmodule
