// Copyright (c) 2015 CERN
// Maciej Suminski <maciej.suminski@cern.ch>
//
// This source code is free software; you can redistribute it
// and/or modify it in source code form under the terms of the GNU
// General Public License as published by the Free Software
// Foundation; either version 2 of the License, or (at your option)
// any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA


// Test for array query functions applied to localparams.

module lparam_query;
localparam const_param = 16'b0001110111001111;

initial begin
    if($left(const_param) !== 15) begin
        $display("FAILED 1");
        $finish();
    end

    if($right(const_param) !== 0) begin
        $display("FAILED 2");
        $finish();
    end

    if($high(const_param) !== 15) begin
        $display("FAILED 3");
        $finish();
    end

    if($low(const_param) !== 0) begin
        $display("FAILED 4");
        $finish();
    end

    if($increment(const_param) !== 1) begin
        $display("FAILED 5");
        $finish();
    end

    if($size(const_param) !== 16) begin
        $display("FAILED 6");
        $finish();
    end

    $display("PASSED");
end
endmodule
