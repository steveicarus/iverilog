module cb();

always begin
  #1;
end

endmodule
