module top;
  initial begin : named_begin
    $display("FAILED");
  end : wrong_name
endmodule
