module tb;
initial $finish(0);
final $display("In final statement.");
endmodule
