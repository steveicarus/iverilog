module test();

logic [1:0] array = new[4];

endmodule
