module a();
endmodule

module test();
a a();
endmodule

module a();
endmodule

module b();
endmodule
