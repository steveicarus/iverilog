// Regression test for GitHub issue #60 part 1 - sized numeric constants
// must have size greater than zero.

module test();

localparam Value = 0'b0;

endmodule
