module top_module();

integer Value1;

parameter Value2 = Value1;

endmodule
