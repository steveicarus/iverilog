// Check a global timeprecision that is too large.
`resetall
timeunit 1ns/10ns;
module gtp_large;
endmodule

