module top;
  parameter value = (1:2:3);
  initial $display(value);
endmodule
