// Check that declarations for dynamic arrays of queues are supported.

module test;

  // Dynamic array of queues
  int q[$][];

endmodule
