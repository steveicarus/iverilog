module top;
  parameter real rpar1 = 1.0;
  parameter real rpar2 = 2.0;
  parameter real rparb = {rpar1, rpar2};
  parameter real rpar = {2.0, 1.0};
endmodule
