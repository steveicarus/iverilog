module test ( input a, input _b_, output A, output b__);
  assign A = a;
  assign b__ = _b_;
endmodule
