module test();

initial
    $display("Error: %m");
endmodule
