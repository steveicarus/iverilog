module top_module();

integer N;

(* attr = N *)
initial $display(N);

endmodule
