// Check that declarations for unpacked arrays of queues are supported.

module test;

  // Unpacked array of queues
  int q[$][10];

endmodule
