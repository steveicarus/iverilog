`define world World
`define test Hello `world

module test;
   initial $display("The `test definition is: `define %s", ``test);
endmodule
