module test;
wire s1;
not(,s1);
not(s1,);
endmodule
