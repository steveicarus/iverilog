// Check that it is an error to declare a non-ANSI task port with implicit
// packed dimensions if it is later redeclared as an integer typed variable.
// Even if the size of the packed dimensions matches that of the size of the
// integer type.

module test;

  task t;
    input [31:0] x;
    integer x;
    $display("FAILED");
  endtask

  initial t(10);

endmodule
