/*
 * Copyright (c) 1999-2000 Stephen Williams (steve@icarus.com)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 */

/*
 * This is derived from pr602.
 */

module main;

   reg [1:0] a [3:0], x;

   integer   i;
   initial begin
      a[0] = 0;
      a[1] = 1;
      a[2] = 2;
      a[3] = 3;

      // The index expressions of this parameter expression
      // should be evaluated to constants.
      $display("a[(1-1)+0] = %b", a[(1-1)+0]);
      $display("a[(2-1)+0] = %b", a[(2-1)+0]);
      x =  a[(1-1)+0];
      if (x !== 2'b00) begin
	 $display("FAILED -- x == %b", x);
	 $finish;
      end

      x =  a[(2-1)+0];
      if (x !== 2'b01) begin
	 $display("FAILED -- x == %b", x);
	 $finish;
      end

      x <=  a[(1-1)+0];
      #1 if (x !== 2'b00) begin
	 $display("FAILED -- x == %b", x);
	 $finish;
      end

      x <=  a[(2-1)+0];
      #1 if (x !== 2'b01) begin
	 $display("FAILED -- x == %b", x);
	 $finish;
      end

      $display("PASSED");
   end // initial begin
endmodule // main
