`define TESTFILE "ivltests/pr3012758.inc"
module top;
`include `TESTFILE
endmodule
