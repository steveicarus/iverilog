`ifndef FOO
`define FOO
`define BAR(x)
`endif

module macro_args();
	macro_args_sub sub();
endmodule
