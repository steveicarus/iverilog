module module_0 (
    id_2,
    id_3,
    id_18,
);
  inout id_18;
  input id_3;
  inout id_2;
  assign id_18 = id_3.id_2;
endmodule
