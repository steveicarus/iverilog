//
// Copyright (c) 1999 Steven Wilson (stevew@home.com)
//
//    This source code is free software; you can redistribute it
//    and/or modify it in source code form under the terms of the GNU
//    General Public License as published by the Free Software
//    Foundation; either version 2 of the License, or (at your option)
//    any later version.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program; if not, write to the Free Software
//    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
//
//  SDW - Validate always #1 disable task_identifier ;

module main ;


reg [3:0] value1 ;

task foo ;
  value1 = #2  1;
endtask

initial
  begin
    value1 = 1'b0;
    #5;
    foo ;
    #4 ;
    if(value1 === 1'b0)
      $display("PASSED");
    else
      $display("FAILED - always3.1.9C always #2 disable foo");
    $finish ;
  end

always #6 disable foo ;

endmodule
