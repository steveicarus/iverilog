module test;
  // For now we just parse these and do not actually do anything with them
  // See section IEEE1800-2012: section 6.9.2
  wire scalared [7:0] scl;
  wire vectored [7:0] vec;

  initial $display("PASSED");
endmodule
