module test;
   initial
     begin
	if(2)
	  $display("PASSED");
	else
	  $display("FAILED");
     end

 endmodule
