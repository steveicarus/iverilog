/*
 * Copyright (c) 2002 Stephen Williams (steve@icarus.com)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 */
module test();

   reg  [7:0]  test;
   wire [7:0]  neg_test = -test;

   initial begin
      for (test = 0 ;  test < 255 ;  test = test + 1) begin
	 #1 if (neg_test !== (-test)) begin
	    $display("FAILED -- %b !== -%b", neg_test, test);
	    $finish;
	 end
      end

      $display("PASSED");
   end

endmodule
