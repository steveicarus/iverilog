module top_module();

integer Value1;

integer Value2 = Value1;

initial $display("PASSED");

endmodule
