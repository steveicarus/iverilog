// Check that declarations for unpacked arrays of dynamic arrays are supported.

module test;

  // Unpacked array of dynamic arrays
  int q[][10];

endmodule
