module top;
  parameter WIDTH = dut.WIDTH;

  test dut();
endmodule

module test;
  parameter WIDTH = 8;
endmodule
