package p1;

endpackage

package p2;

logic x;

endpackage

module m;

initial $dumpvars;

endmodule
