module top;
  buf sclbuf0();
endmodule
