//
// Copyright (c) 1999 Steven Wilson (stevew@home.com)
//
//    This source code is free software; you can redistribute it
//    and/or modify it in source code form under the terms of the GNU
//    General Public License as published by the Free Software
//    Foundation; either version 2 of the License, or (at your option)
//    any later version.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program; if not, write to the Free Software
//    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
//
//  SDW - Validate 3 way fork. Bug report 228.

module test;

reg a,b,c;
reg error;


initial
  begin
    error = 0;
    fork
      a = 1;
      b = 0;
      c = 1;
    join

  if(a !== 1)
     begin
       $display("FAILED - a not set to 1");
       error = 1;
     end
  if(b !== 0)
     begin
       $display("FAILED - b not set to 0");
       error = 1;
     end
  if(c !== 1)
     begin
       $display("FAILED - c not set to 1");
       error = 1;
     end
  if(error == 0)
    $display("PASSED");

  end

endmodule
