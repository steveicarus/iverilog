// pr1960548

module test;
   initial
     $display("B`x");
endmodule
