// Check a missing global time precision.
`resetall
timeunit 1ns;
module no_gtp;
endmodule
