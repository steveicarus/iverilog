module test();

`define MACRO 1
`define MACRO 1
`define MACRO 2
`undef MACRO
`define MACRO 1

endmodule
