/*
 * Copyright (c) 2002 Stephen Williams (steve@icarus.com)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 */

/*
 */
`timescale 1ns / 1ns

module main;

   initial begin
      #3 $display("$time = %t (unformatted)", $time);
      $timeformat(-6, 6, "ns", 12);
      $display("$time = %t (-6,6)", $time);
      $timeformat(-6, 1, "ns", 12);
      $display("$time = %t (-6,1)", $time);
   end


endmodule // main
