module test();

reg [7:0] ival = $signed(1.0);

endmodule
