module if_fail_test();

`ifdef
`ifndef
`elsif
`else
`endif

  initial $display("FAILED");

endmodule
