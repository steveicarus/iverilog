module t;
  final $display("Final in %m");
endmodule

module t2;
  final $display("Final in %m");
endmodule
