// Check that declarations for dynamic arrays of unpacked arrays are supported.

module test;

  // Dynamic array of unpacked arrays
  int q[10][];

endmodule
