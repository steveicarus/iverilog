module top;
  reg var;

  always if (var);
endmodule
