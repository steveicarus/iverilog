module top;
  initial begin : named_begin
    $display("PASSED");
  end : named_begin
endmodule
