module test();

wire real r;

assign r = 1.0;
assign r = 2.0;

endmodule
