module top;
  specify
    specparam s_int = -1;
    specparam s_real = -1.0;
 endspecify
endmodule
