module test();

wire bit [7:0] b;

assign b = 8'h11;
assign b = 8'h22;

endmodule
