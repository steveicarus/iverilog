// Check that declarations for queues of dynamic arrays are supported.

module test;

  // Queue of dynamic arrays
  int q[][$];

endmodule
