(* foo, bar=1 *) (* baz=1 *) module foo;
  initial $display("PASSED");
endmodule
