module test();

reg illegal[0];

endmodule
