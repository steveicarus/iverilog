module test;

initial $display("FAILED");

endmodule
