// Check that declarations for queues of queues are supported.

module test;

  // Queue of queues
  int q[$][$];

endmodule
