module top;
  initial begin
    logic [7:0] data;
    logic [3:0] tmp;
  end

  initial begin
    logic [3:0] nib;
    $display("PASSED");
  end
endmodule
