//
// Copyright (c) 2000 Paul Campbell (paul@verifarm.com)
//
//    This source code is free software; you can redistribute it
//    and/or modify it in source code form under the terms of the GNU
//    General Public License as published by the Free Software
//    Foundation; either version 2 of the License, or (at your option)
//    any later version.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program; if not, write to the Free Software
//    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
//
module compl1000;
	reg	[158:143]r0;
	reg	[128:104]r1;
	reg	[200:173]r2;
	reg	[165:162]r3;
	reg	[150:129]r4;
	reg	[123:93]r5;
	reg	[55:54]r6;
	reg	[24:3]r7;
	reg	[109:93]r8;
	reg	[30:14]r9;
	reg	[184:174]r10;
	reg	[59:30]r11;
	reg	[153:124]r12;
	reg	[248:221]r13;
	reg	[258:250]r14;
	reg	[158:147]r15;
	reg	[54:48]r16;
	reg	[159:136]r17;
	reg	[214:187]r18;
	reg	[60:29]r19;
	reg	[71:71]r20;
	reg	[177:169]r21;
	reg	[219:205]r22;
	reg	[24:21]r23;
	reg	[153:141]r24;
	reg	[85:54]r25;
	reg	[227:202]r26;
	reg	[251:237]r27;
	reg	[98:73]r28;
	reg	[24:0]r29;
	reg	[166:135]r30;
	reg	[184:183]r31;
	reg	[219:189]r32;
	reg	[81:54]r33;
	reg	[164:148]r34;
	reg	[170:158]r35;
	reg	[171:168]r36;
	reg	[255:226]r37;
	reg	[197:191]r38;
	reg	[113:105]r39;
	reg	[221:198]r40;
	reg	[135:104]r41;
	reg	[153:143]r42;
	reg	[281:253]r43;
	reg	[101:76]r44;
	reg	[24:12]r45;
	reg	[217:203]r46;
	reg	[244:218]r47;
	reg	[128:111]r48;
	reg	[136:107]r49;
	reg	[260:242]r50;
	reg	[157:156]r51;
	reg	[242:220]r52;
	reg	[278:255]r53;
	reg	[196:194]r54;
	reg	[148:121]r55;
	reg	[71:63]r56;
	reg	[166:157]r57;
	reg	[200:180]r58;
	reg	[230:199]r59;
	reg	[212:191]r60;
	reg	[264:248]r61;
	reg	[136:124]r62;
	reg	[131:117]r63;
	reg	[148:126]r64;
	reg	[51:30]r65;
	reg	[166:140]r66;
	reg	[166:143]r67;
	reg	[44:27]r68;
	reg	[259:248]r69;
	reg	[167:143]r70;
	reg	[210:189]r71;
	reg	[73:50]r72;
	reg	[225:205]r73;
	reg	[255:240]r74;
	reg	[208:194]r75;
	reg	[222:217]r76;
	reg	[217:189]r77;
	reg	[100:83]r78;
	reg	[275:255]r79;
	reg	[39:34]r80;
	reg	[98:72]r81;
	reg	[55:25]r82;
	reg	[246:240]r83;
	reg	[170:157]r84;
	reg	[218:198]r85;
	reg	[225:223]r86;
	reg	[186:172]r87;
	reg	[241:213]r88;
	reg	[263:238]r89;
	reg	[272:253]r90;
	reg	[105:103]r91;
	reg	[211:209]r92;
	reg	[89:82]r93;
	reg	[30:9]r94;
	reg	[246:241]r95;
	reg	[170:147]r96;
	reg	[229:224]r97;
	reg	[107:83]r98;
	reg	[60:54]r99;
	reg	[154:154]r100;
	reg	[105:97]r101;
	reg	[127:104]r102;
	reg	[219:190]r103;
	reg	[114:98]r104;
	reg	[267:251]r105;
	reg	[169:145]r106;
	reg	[64:45]r107;
	reg	[227:224]r108;
	reg	[186:176]r109;
	reg	[101:84]r110;
	reg	[219:194]r111;
	reg	[11:9]r112;
	reg	[236:222]r113;
	reg	[271:240]r114;
	reg	[232:218]r115;
	reg	[78:74]r116;
	reg	[191:191]r117;
	reg	[242:227]r118;
	reg	[135:108]r119;
	reg	[24:15]r120;
	reg	[250:233]r121;
	reg	[125:102]r122;
	reg	[165:140]r123;
	reg	[63:63]r124;
	reg	[235:206]r125;
	reg	[264:237]r126;
	reg	[241:234]r127;
	reg	[188:188]r128;
	reg	[71:59]r129;
	reg	[181:170]r130;
	reg	[106:83]r131;
	reg	[245:229]r132;
	reg	[239:219]r133;
	reg	[10:8]r134;
	reg	[45:45]r135;
	reg	[23:22]r136;
	reg	[197:178]r137;
	reg	[57:50]r138;
	reg	[264:253]r139;
	reg	[53:36]r140;
	reg	[187:164]r141;
	reg	[153:140]r142;
	reg	[235:226]r143;
	reg	[236:228]r144;
	reg	[262:238]r145;
	reg	[76:55]r146;
	reg	[49:25]r147;
	reg	[191:163]r148;
	reg	[197:170]r149;
	reg	[151:143]r150;
	reg	[126:122]r151;
	reg	[188:173]r152;
	reg	[93:78]r153;
	reg	[175:175]r154;
	reg	[249:247]r155;
	reg	[214:200]r156;
	reg	[60:43]r157;
	reg	[263:233]r158;
	reg	[54:34]r159;
	reg	[202:184]r160;
	reg	[250:240]r161;
	reg	[99:80]r162;
	reg	[175:165]r163;
	reg	[189:188]r164;
	reg	[52:38]r165;
	reg	[74:48]r166;
	reg	[232:202]r167;
	reg	[24:13]r168;
	reg	[209:180]r169;
	reg	[173:147]r170;
	reg	[264:243]r171;
	reg	[115:99]r172;
	reg	[94:91]r173;
	reg	[195:188]r174;
	reg	[36:33]r175;
	reg	[136:114]r176;
	reg	[82:56]r177;
	reg	[204:173]r178;
	reg	[116:111]r179;
	reg	[124:103]r180;
	reg	[76:71]r181;
	reg	[178:163]r182;
	reg	[156:149]r183;
	reg	[124:110]r184;
	reg	[240:220]r185;
	reg	[164:151]r186;
	reg	[133:104]r187;
	reg	[59:46]r188;
	reg	[47:42]r189;
	reg	[219:189]r190;
	reg	[99:87]r191;
	reg	[86:73]r192;
	reg	[222:191]r193;
	reg	[23:7]r194;
	reg	[239:238]r195;
	reg	[240:222]r196;
	reg	[27:4]r197;
	reg	[191:160]r198;
	reg	[106:84]r199;
	reg	[22:8]r200;
	reg	[204:191]r201;
	reg	[133:115]r202;
	reg	[225:207]r203;
	reg	[126:95]r204;
	reg	[161:147]r205;
	reg	[193:164]r206;
	reg	[69:61]r207;
	reg	[130:116]r208;
	reg	[142:124]r209;
	reg	[50:20]r210;
	reg	[175:154]r211;
	reg	[102:87]r212;
	reg	[114:85]r213;
	reg	[225:223]r214;
	reg	[131:127]r215;
	reg	[24:19]r216;
	reg	[84:84]r217;
	reg	[223:223]r218;
	reg	[171:159]r219;
	reg	[76:47]r220;
	reg	[162:139]r221;
	reg	[67:41]r222;
	reg	[88:74]r223;
	reg	[60:44]r224;
	reg	[114:104]r225;
	reg	[142:141]r226;
	reg	[262:236]r227;
	reg	[16:12]r228;
	reg	[66:51]r229;
	reg	[40:24]r230;
	reg	[150:141]r231;
	reg	[209:199]r232;
	reg	[152:148]r233;
	reg	[162:147]r234;
	reg	[82:80]r235;
	reg	[245:214]r236;
	reg	[35:12]r237;
	reg	[18:3]r238;
	reg	[270:246]r239;
	reg	[183:170]r240;
	reg	[122:121]r241;
	reg	[60:42]r242;
	reg	[99:91]r243;
	reg	[61:51]r244;
	reg	[154:150]r245;
	reg	[5:3]r246;
	reg	[275:246]r247;
	reg	[113:92]r248;
	reg	[136:118]r249;
	reg	[94:71]r250;
	reg	[104:91]r251;
	reg	[169:139]r252;
	reg	[22:14]r253;
	reg	[255:236]r254;
	reg	[213:186]r255;
	initial begin
		r0 = 32'h3d24;
		r1 = 32'h70fd;
		r2 = 32'h47aa;
		r3 = 32'h39ed;
		r4 = 32'h2ca3;
		r5 = 32'he68;
		r6 = 32'h1160;
		r7 = 32'h5636;
		r8 = 32'h2305;
		r9 = 32'h1257;
		r10 = 32'h4e74;
		r11 = 32'h3835;
		r12 = 32'h3857;
		r13 = 32'h3f6f;
		r14 = 32'h7b33;
		r15 = 32'h2f37;
		r16 = 32'h10a;
		r17 = 32'h6cff;
		r18 = 32'h3f3;
		r19 = 32'h70e2;
		r20 = 32'h4cb3;
		r21 = 32'h510;
		r22 = 32'h1837;
		r23 = 32'h425;
		r24 = 32'h1488;
		r25 = 32'h5731;
		r26 = 32'h1388;
		r27 = 32'h6ee0;
		r28 = 32'h559b;
		r29 = 32'h4bff;
		r30 = 32'h180e;
		r31 = 32'h1252;
		r32 = 32'h52d4;
		r33 = 32'h4576;
		r34 = 32'h36f1;
		r35 = 32'h6246;
		r36 = 32'h7aaf;
		r37 = 32'h37fb;
		r38 = 32'h4272;
		r39 = 32'h62fd;
		r40 = 32'h6cbb;
		r41 = 32'h4825;
		r42 = 32'h25c7;
		r43 = 32'h19da;
		r44 = 32'h5ace;
		r45 = 32'h794f;
		r46 = 32'h5ebb;
		r47 = 32'h5cd0;
		r48 = 32'h4209;
		r49 = 32'h38de;
		r50 = 32'h7502;
		r51 = 32'h2c8c;
		r52 = 32'h378f;
		r53 = 32'h5252;
		r54 = 32'hb5d;
		r55 = 32'h561;
		r56 = 32'h4504;
		r57 = 32'h180f;
		r58 = 32'h6672;
		r59 = 32'h52f7;
		r60 = 32'h10c7;
		r61 = 32'h4ce9;
		r62 = 32'h569;
		r63 = 32'h72b3;
		r64 = 32'h4df0;
		r65 = 32'h1a72;
		r66 = 32'h2846;
		r67 = 32'h70e5;
		r68 = 32'h3008;
		r69 = 32'h2003;
		r70 = 32'h6009;
		r71 = 32'h6cb5;
		r72 = 32'h5e8b;
		r73 = 32'h668b;
		r74 = 32'h487;
		r75 = 32'h4eca;
		r76 = 32'h241e;
		r77 = 32'h451a;
		r78 = 32'h2c06;
		r79 = 32'h3ebf;
		r80 = 32'h5590;
		r81 = 32'h22c;
		r82 = 32'h9b;
		r83 = 32'h347;
		r84 = 32'h2c92;
		r85 = 32'h3db6;
		r86 = 32'hf44;
		r87 = 32'h391a;
		r88 = 32'h1237;
		r89 = 32'h6ff2;
		r90 = 32'h6cc5;
		r91 = 32'hca7;
		r92 = 32'h152a;
		r93 = 32'h8eb;
		r94 = 32'h4c43;
		r95 = 32'h6277;
		r96 = 32'h7b1;
		r97 = 32'h7cc8;
		r98 = 32'h63a2;
		r99 = 32'h1a62;
		r100 = 32'h165;
		r101 = 32'h48d8;
		r102 = 32'h399e;
		r103 = 32'h5975;
		r104 = 32'h40ae;
		r105 = 32'h3d61;
		r106 = 32'h39ab;
		r107 = 32'h69f;
		r108 = 32'h2801;
		r109 = 32'h1828;
		r110 = 32'h298d;
		r111 = 32'h661e;
		r112 = 32'h52d9;
		r113 = 32'h3bc0;
		r114 = 32'h5cb7;
		r115 = 32'h7fac;
		r116 = 32'h7e76;
		r117 = 32'hf93;
		r118 = 32'h4165;
		r119 = 32'h3b68;
		r120 = 32'h4258;
		r121 = 32'h54b2;
		r122 = 32'h2378;
		r123 = 32'h6186;
		r124 = 32'h547a;
		r125 = 32'h7b5c;
		r126 = 32'h4115;
		r127 = 32'h68b6;
		r128 = 32'h554f;
		r129 = 32'h4550;
		r130 = 32'hcfc;
		r131 = 32'h3f55;
		r132 = 32'h5f7d;
		r133 = 32'h40d2;
		r134 = 32'h3aa8;
		r135 = 32'h7b56;
		r136 = 32'h575c;
		r137 = 32'h687f;
		r138 = 32'h702c;
		r139 = 32'h1cee;
		r140 = 32'h362d;
		r141 = 32'h73d2;
		r142 = 32'h39c8;
		r143 = 32'h5003;
		r144 = 32'h4d1a;
		r145 = 32'h2472;
		r146 = 32'h1b4e;
		r147 = 32'h5852;
		r148 = 32'h3bf2;
		r149 = 32'h1c41;
		r150 = 32'h5b37;
		r151 = 32'h1462;
		r152 = 32'h17a1;
		r153 = 32'h825;
		r154 = 32'h6384;
		r155 = 32'h432c;
		r156 = 32'h7c70;
		r157 = 32'h2b94;
		r158 = 32'h5456;
		r159 = 32'h7887;
		r160 = 32'h802;
		r161 = 32'h18e2;
		r162 = 32'h244c;
		r163 = 32'h6c55;
		r164 = 32'h770a;
		r165 = 32'h224a;
		r166 = 32'h6aa0;
		r167 = 32'h1070;
		r168 = 32'h62cd;
		r169 = 32'h4fbe;
		r170 = 32'h2f01;
		r171 = 32'h1952;
		r172 = 32'h5a5b;
		r173 = 32'h656e;
		r174 = 32'h5b2e;
		r175 = 32'h6586;
		r176 = 32'h538d;
		r177 = 32'h471a;
		r178 = 32'h2a57;
		r179 = 32'h6fd2;
		r180 = 32'h2fbd;
		r181 = 32'h4418;
		r182 = 32'h3233;
		r183 = 32'h3821;
		r184 = 32'h5048;
		r185 = 32'h1824;
		r186 = 32'h61e0;
		r187 = 32'h4f33;
		r188 = 32'h76c5;
		r189 = 32'h2ceb;
		r190 = 32'h127f;
		r191 = 32'h7103;
		r192 = 32'h6d02;
		r193 = 32'h6856;
		r194 = 32'h58b;
		r195 = 32'h59fb;
		r196 = 32'h30c3;
		r197 = 32'h1397;
		r198 = 32'h6cfd;
		r199 = 32'h42da;
		r200 = 32'h1f39;
		r201 = 32'h26f4;
		r202 = 32'h5922;
		r203 = 32'h2f61;
		r204 = 32'h5c44;
		r205 = 32'h656;
		r206 = 32'h2837;
		r207 = 32'h7bc1;
		r208 = 32'h7168;
		r209 = 32'h7a91;
		r210 = 32'h53ca;
		r211 = 32'h54c4;
		r212 = 32'h6091;
		r213 = 32'h7371;
		r214 = 32'h37d0;
		r215 = 32'h6bd;
		r216 = 32'h2687;
		r217 = 32'h5e88;
		r218 = 32'h2f85;
		r219 = 32'h4f31;
		r220 = 32'h692f;
		r221 = 32'h1eba;
		r222 = 32'h2407;
		r223 = 32'h1d42;
		r224 = 32'h4d87;
		r225 = 32'h7085;
		r226 = 32'h68b1;
		r227 = 32'h6cdf;
		r228 = 32'h315f;
		r229 = 32'h4711;
		r230 = 32'h138;
		r231 = 32'h28ad;
		r232 = 32'h44d8;
		r233 = 32'h6dfb;
		r234 = 32'h2d88;
		r235 = 32'h3eb4;
		r236 = 32'h3f9e;
		r237 = 32'h7be1;
		r238 = 32'h575c;
		r239 = 32'h53ca;
		r240 = 32'h2de5;
		r241 = 32'h61ad;
		r242 = 32'h3d9f;
		r243 = 32'h41c0;
		r244 = 32'h1124;
		r245 = 32'h22a2;
		r246 = 32'h7986;
		r247 = 32'h4c4e;
		r248 = 32'h5094;
		r249 = 32'h128;
		r250 = 32'h396a;
		r251 = 32'h38be;
		r252 = 32'h3567;
		r253 = 32'h2c57;
		r254 = 32'h4d66;
		r255 = 32'h345b;
		#10; r201 = $stime;
		#10; r153 =  ( ~ ( r189));
		#10; r200 = (3'h7 !== r2);
		#10; r186 = r155;
		#10; r208 = (((((( ( + ( (((16'h46d9 || r190) - $time) > (r127 >= (2'h0 !== r81))))) ||  ( | ( r150))) > r11) !== ((20'h617c *  ( & ( r207))) > (r158 && (31'h6f3f - 19'h3eb3)))) * 17'h5321) - 25'h116f) ^ ((((($stime === r219) <= ($stime | (r43 < ((($stime ^ (( ( & ( ( ( & ( 26'h3af4)) |  ( | ( 12'h8c7))))) && (r97 | 7'h3)) && 17'h7a8a)) == 9'h84) + ((18'h7e64 >= r240) >= r111))))) ^ 8'ha9) ^  ( - ( r15))) & (( ( & ( $time)) == r235) >= (( ( | ( r90)) || (r56 & r182)) !== r72))));
		#10; r175 = (($time / ((15'h7f3d === ( ( & ( r1)) == r2)) >= ((9'h78 % ( ( ^ (  ( - ( (r164 & (2'h2 >= (((((6'h1f == 28'h4032) /  ( | ( 16'h5821))) | 28'h7b43) >= (r191 & $stime)) <  ( + ( ((2'h3 % (12'hf20 - 16'h2734)) ?  ( + ( (16'h1317 && 31'h16ee))) : (r137 < (6'h27 >= 3'h2)))))))))))) & ((( ( - ( (r169 ? ((r155 != 31'h60f0) >= ((r166 % (15'h587f - 30'h5197)) < r187)) : (((23'h220b <= 20'h46a) & (29'h584 > (10'h17 - 19'h53b7))) !=  ( & (  ( | ( (9'h1d0 <= 2'h0))))))))) ? r92 : ((($time <= 27'h6600) < (5'h13 ^ r99)) <=  ( ! ( (((17'h2640 ? 2'h1 : r189) > $time) >= r248))))) ? (3'h2 - (9'h97 ==  ( ^ ( 4'h5)))) : ((1'h0 ? ( ( ! ( r34)) && ((r61 >= r73) == ((r184 === (19'h2c6c != 19'h34df)) |  ( ~ ( r72))))) : 19'h64ff) >= (( ( ! ( (r24 !== ((7'h2b >= 1'h1) &&  ( ~ ( 4'he)))))) <=  ( ^ ( r86))) / 12'hff3))) % (r35 <  ( - ( 13'h8b9)))))) && r67))) - (((8'h12 !== (14'h2d97 <= ((r183 !== (((((r19 | r178) | (32'h743d != (r199 > ((28'h6bbb - 9'hc1) /  ( + ( 18'h25d4)))))) | r255) < ( ( | ( (r12 | ((r255 % (30'h5e7b >= 11'h753)) < ( ( ~ ( 29'hc71)) || (20'h1ffc <= 17'h7cc5)))))) !== ((r181 * (((11'h18f || 17'h7265) ? 29'h485f : 4'he) == ( ( ~ ( 14'h1c84)) + 23'h298c))) || (((20'h79b3 ? (25'h1681 * 4'h9) : (12'ha6e * 26'h3ed1)) <= (r84 | (1'h1 % 2'h3))) ^ (r0 < ( ( ! ( 10'h336)) % (10'h149 / 3'h4))))))) || (r184 <= 26'h55e8))) ? 5'h17 :  ( & ( (1'h0 >= r248)))))) + r191) | r65));
		#10; r28 = ( ( ! ( ($time <= r162))) !== r91);
		#10; r125 = ($stime ===  ( - ( r231)));
		#10; r237 = r93;
		#10; r150 = (( ( - ( r183)) &  ( ~ ( (23'h3dd8 === $time)))) > r75);
		#10; r59 = (23'h7ddf * $stime);
		#10; r157 = (3'h4 + (r27 |  ( ^ ( (r175 ^ 8'h7b)))));
		#10; r65 = r109;
		#10; r241 = r88;
		#10; r96 = 7'h62;
		#10; r229 = (r248 + (r37 >= $time));
		#10; r112 = r160;
		#10; r73 = 26'h5f00;
		#10; r72 = r17;
		#10; r2 = ( ( | ( (r124 + (( ( | ( (7'hf && (r196 ? r84 : ( ( & ( r51)) / r215))))) <= r7) <=  ( | ( (r250 + ((20'h6268 % r214) / r19)))))))) * ( ( ! ( ((r249 % ($stime && (r140 *  ( - ( ((r104 / 4'h4) <= (( ( + ( r250)) -  ( | ( r68))) &  ( ~ ( $time))))))))) || (r96 > (23'h4f58 < r185))))) !== 27'h5720));
		#10; r66 = r133;
		#10; r199 =  ( & ( (r2 %  ( ^ (  ( - (  ( - ( r20)))))))));
		#10; r47 = r109;
		#10; r55 = (r96 / (r204 |  ( + ( (((14'h519 / ((32'h2b24 ? ( ( | (  ( ^ ( r184)))) * (r123 < r123)) : ((((((r37 - (5'h13 == 10'h211)) ==  ( ! ( $time))) * 19'h76aa) >= ( ( | ( r211)) != r116)) ^  ( + ( 10'h25c))) ? (31'h68d3 !== (28'h6b7 ? ((($stime ||  ( + ( 25'h7c9a))) | (r74 ===  ( & ( 31'h28e9)))) %  ( + ( ((1'h0 && 28'h6335) |  ( - ( 13'h130c)))))) : 1'h0)) : ((r115 ||  ( | ( ( ( ~ ( r133)) && ((23'h30d3 ^ 32'h4295) % (18'h417d >= 22'h51c3)))))) && (((23'h7803 != ( ( ! ( 14'h1906)) ^ (19'h837 > 2'h2))) * (r198 <= (23'h1ee0 <= r55))) >= $stime)))) < ( ( ^ ( ((16'h5ded | (r217 / 17'h171e)) || 1'h0))) > r250))) < (8'h89 && (r15 |  ( - ( r224))))) !== (((r244 === (((r229 <= 28'h441b) - ( ( | ( ((r244 - ((29'h24d7 != 17'h334f) == (8'h9f ^ 32'h3180))) ^  ( ^ ( (r238 * (21'h5f35 / 20'h5115))))))) * ( ( + (  ( - (  ( ~ ( (19'h79a9 ^ 24'h5d6a))))))) % r113))) > (((((r92 * (r232 * (22'h261f <= 14'h2bc3))) & (((20'h309a & 22'h7de2) && r181) < ((19'h7534 | 29'h18ae) > r188))) == ((((13'h46f && 25'h1d09) % r161) -  ( ^ ( 30'h7cd8))) +  ( - ( ((22'h6d8b || 29'h3b) ^ (21'h24f3 > 8'h7f)))))) | (r59 && (r191 >= ( ( & ( (12'h473 & 7'h69))) <= ((30'h162e !== 27'h1a0d) | 18'h5c9a))))) & (r182 - (( ( ~ ( (23'h70cb * (24'h246d > 2'h1)))) - (( ( & ( 26'h6e6c)) == 28'h21af) !== 8'h6f)) % (4'h4 >= r168)))))) != (( ( ~ ( r31)) && ( ( + ( r130)) / r96)) > 19'h1be5)) /  ( ~ (  ( + ( ( ( ! ( (((r154 ? (r253 !==  ( | ( (1'h0 % 22'h7fd4)))) : ((r133 > (29'h70f ? 6'h3a : 19'hff4)) === 26'h9dd)) <= r109) != 4'h2))) *  ( & ( 4'h4)))))))))))));
		#10; r70 = r113;
		#10; r111 =  ( ! ( ( ( ^ (  ( - (  ( | (  ( | ( ((r207 * ((((r224 !== (15'h2f78 < 32'h5844)) > (r246 ===  ( + (  ( ! ( r150)))))) >= r24) && 2'h1)) * r208))))))))) || ( ( ^ ( ((((r144 % r39) <  ( - ( ((9'h103 + ( ( & (  ( ~ ( (r176 || (2'h1 ^ 3'h1)))))) ? $stime : r132)) ^  ( + ( (27'h3a07 ? ( ( ^ ( r12)) && ( ( & ( r164)) -  ( + ( (2'h0 > 29'h1ec3))))) : r114))))))) && r126) && ((15'h4051 !== (r0 >= 27'h7733)) ^ (((22'h3da3 | ( ( & (  ( ^ ( r90)))) & 2'h1)) / 2'h1) === (r51 % r189)))))) !== (r252 == 4'h5)))));
		#10; r162 = 6'h25;
		#10; r183 = ( ( - ( (r110 ?  ( ^ ( ( ( + ( ((26'h7b30 != 7'h4c) - r124))) * $time))) :  ( + ( (r178 * r22)))))) ^ ((r155 && r52) < (r118 ^ ( ( | ( ( ( ! ( (24'h35fc ^ ((( ( & ( ((r53 - r49) >= 5'ha))) ? r251 : r162) <= 21'h5575) ? (r163 != (( ( ~ ( r203)) - r130) + r153)) : r97)))) == (((r154 |  ( ! ( (r105 | r241)))) !== ((18'h6bbe +  ( ^ ( (r193 !==  ( ^ ( r26)))))) == 6'h1d)) - ((((((((11'h11f || 7'h25) ? r117 : (3'h4 > 19'h2c65)) + ((29'h1842 | 18'h1c77) +  ( | ( 13'h19b)))) == $stime) != 11'h491) - 18'h69a8) & (((r206 ?  ( - ( (30'hd83 ^ (30'h7ac6 | 2'h2)))) : (((10'h9d && 32'h5721) === $time) !== (r190 === (9'hd9 / 27'h2d)))) && (r232 || (r76 >  ( + ( 25'hd8b))))) < $stime)) == r191))))) + $time))));
		#10; r30 = r66;
		#10; r60 = (22'h3eec ^ (11'h1dd ^ 9'h113));
		#10; r229 =  ( ~ ( 5'hc));
		#10; r180 =  ( ^ (  ( & ( r127))));
		#10; r30 = r124;
		#10; r149 =  ( - ( (30'h743 === ((((((13'hc2 * (( ( & ( 30'h12da)) + 26'h7fc3) + ($stime ? ( ( ~ ( 27'h75f6)) | (r62 !==  ( - ( 21'h3b14)))) : r238))) !== (r248 == 30'h7a43)) || 22'hfbe) * $stime) ? r240 : r4) >= (12'hd38 ^ (r147 + ((r36 - 23'h1ed1) ? ((r123 >= ( ( ~ ( (( ( + (  ( ~ ( (15'h32ce / 32'h6ae6))))) | 12'hf22) > $stime))) ? (((r200 == ($stime && r86)) >= (( ( & ( (1'h0 <= 22'h4156))) != 2'h3) === ((r118 && r106) * r249))) || 16'h629a) : (28'h6bec !== r65))) % ((21'h5864 * 2'h0) % $time)) : ((( ( & (  ( ~ (  ( ~ ( (((17'h19fd != 2'h1) > (23'h4f5d & 26'h14e6)) >=  ( & ( r236))))))))) === ( ( ^ ( ((r146 && ( ( + ( 26'h40d8)) % (11'h5ba ? 16'h7254 : 32'h7877))) != 22'h3cba))) !== ( ( - (  ( ! ( r162)))) / 2'h3))) !=  ( ^ ( (r135 &  ( ~ ( (((26'hc01 !== r252) || ((4'hd | 8'h62) >  ( & ( 16'h4d14)))) == 18'h6094))))))) & (( ( ~ ( r147)) > r72) !== 13'h1f75)))))))));
		#10; r173 = 5'h0;
		#10; r103 = $time;
		#10; r239 = $time;
		#10; r23 = r22;
		#10; r77 = ((13'h16b3 ==  ( & ( r9))) /  ( - ( ($time && 5'h1c))));
		#10; r132 = ((r22 >= (r212 ^ (((($stime === ((r241 % (( ( | ( ($time % ((11'h4b7 && 2'h3) >=  ( ! ( 32'h71f5)))))) - $stime) ? (r98 && 2'h3) :  ( ^ ( (21'h384f === 27'h85))))) <=  ( ! ( (20'h4d8 <= $time))))) !== (r147 == (r51 / r226))) | r15) / r114))) ? r208 : (( ( ~ (  ( + ( $stime)))) != r7) == ( ( - (  ( ! ( ( ( - ( ( ( & ( ((( ( ~ ( 22'h2cd1)) != (((14'h176d <= 29'h32ef) + (16'h23d1 != 2'h1)) * ((1'h0 ^ 14'hf5b) + r98))) || r212) === (r154 ? 5'h4 : ((((6'h18 !== 4'h7) / (27'h2c4d & 14'h1ea)) >  ( | ( $time))) > (( ( + ( 22'h2996)) !== 32'h70cf) && (r135 - r79))))))) | (r98 / r221)))) +  ( ^ ( (r198 !== (9'h10d === 7'h11))))))))) -  ( ~ ( 30'h1aa4)))));
		#10; r43 = (28'h3e31 !=  ( - ( ((r204 ?  ( ~ ( r214)) : r7) && 16'h2745))));
		#10; r161 = ($stime % (( ( | ( (r185 %  ( ^ ( r104))))) % ($time * (((r170 | 17'h229d) ? ((($stime >= (23'h16aa & (r64 != ((r100 & (r61 | $stime)) === r136)))) === 27'h349d) ? ((( ( & ( 4'h8)) ?  ( + ( r122)) :  ( ! (  ( ^ ( r70))))) >  ( ~ ( r159))) + r79) : (7'h72 ^ (r55 /  ( + (  ( | (  ( ^ ( ( ( ~ ( (23'h7fda + 10'h17))) *  ( - ( r1)))))))))))) :  ( ! ( ( ( - ( $stime)) %  ( ~ ( 5'h2)))))) >= ( ( ^ ( r226)) * r107)))) <= 31'h78c1));
		#10; r132 = ((1'h0 === r227) != 24'h6058);
		#10; r128 = 3'h1;
		#10; r15 = 19'h5239;
		#10; r17 = 15'ha01;
		#10; r77 = ((r242 === r221) * (r179 !== r249));
		#10; r87 = (32'h57ec | r63);
		#10; r116 = r136;
		#10; r20 = r148;
		#10; r53 = 30'h6650;
		#10; r140 = r198;
		#10; r246 = ($stime / ( ( | ( $stime)) / ( ( ! (  ( + ( r215)))) & 20'h3e0e)));
		#10; r69 = r246;
		#10; r172 = r163;
		#10; r94 = r157;
		#10; r107 = $stime;
		#10; r74 =  ( + (  ( - ( $time))));
		#10; r130 = r195;
		#10; r197 = (29'ha48 > ((((r121 ^ r165) <= r124) & r226) ^ ((((((r79 * ( ( ~ ( (4'h7 !=  ( ~ ( r188))))) ^ r70)) & ( ( & ( ((r140 - ( ( ! ( ((32'h6c24 >= 7'h2d) == (2'h1 || 32'h1866)))) || 29'h16f1)) > (2'h1 ||  ( + ( ($stime == (r68 | 11'h34b)))))))) == r193)) !== r211) | r227) % (r16 == (r10 && (r229 / 4'hc)))) + (r242 ^ r117))));
		#10; r130 = (20'h23ae | 18'h14b8);
		#10; r136 = 9'h20;
		#10; r249 = 15'h1805;
		#10; r224 = 1'h0;
		#10; r47 = r200;
		#10; r153 = 21'h2587;
		#10; r137 = 29'h4926;
		#10; r241 =  ( | ( (r228 ? ((((27'h60f7 <  ( ^ ( ( ( ^ (  ( - ( (r82 / 8'hb9))))) & ( ( ^ ( r124)) >= (r222 ^ (($stime ^  ( & (  ( ! ( 8'h30))))) * r146))))))) == r4) | ($time % (1'h0 /  ( | ( (( ( | (  ( ^ ( ((( ( ^ ( 29'h3ca3)) / (8'h37 == 26'h3dbc)) + ((30'h160b >= 23'h7433) ^ r114)) >= (18'h2332 ? (20'h14e1 / (18'h1626 && 28'h64b1)) : r88)))))) < r219) ^ ( ( - (  ( & (  ( + ( ( ( ! ( (25'h7e80 | 5'h14))) >  ( - ( (16'h12d2 || 9'h1c2)))))))))) ? $time : $stime))))))) !== r104) : ((((r252 || r121) | ((6'h37 == (((17'h697e === r43) + (18'h44f4 % 5'h1a)) ? r117 : r30)) < $stime)) + ((((r167 ?  ( | ( (r87 +  ( ! ( (19'h6a46 < r109)))))) :  ( ! ( 16'hb75))) == 32'h4122) | r99) / (((15'h25b8 ===  ( ^ ( r158))) == ( ( ~ ( 23'h693a)) -  ( | (  ( ^ ( r249)))))) / (r168 ? ( ( ^ ( r95)) - $time) : r204)))) * (r139 !== 24'h3813)))));
		#10; r166 = ( ( - ( ((r111 === r215) && r112))) | ((((($stime != r97) / ((22'h6297 != (((20'h58b | (r76 ? $time : (r57 > (( ( - ( 22'h52e5)) - (14'h105e === 4'hc)) ^  ( & ( (28'h7a38 || 14'h3a92))))))) | (23'h2ee7 / (r70 + r159))) > 17'h862)) >= (24'h4bd6 > $stime))) < (((((22'h38cf * r181) -  ( + ( (r36 == r49)))) !== 18'h15e4) & r185) ^  ( ^ ( 19'h2b9c)))) ==  ( & ( r150))) ==  ( & ( r137))));
		#10; r236 = ( ( + ( ((((((r148 || ( ( ~ (  ( - (  ( ~ ( r254)))))) != (6'h20 <= r133))) > 26'h163c) !==  ( & ( (($time === r13) != 15'h637b)))) === 24'h7118) <  ( + ( r42))) / r251))) ? (r43 % (6'h2 ===  ( + ( r209)))) : ($stime ==  ( + ( r82))));
		#10; r35 = 32'h194c;
		#10; r242 = 12'h485;
		#10; r163 = r152;
		#10; r143 = (r53 >= ((r240 || 4'h8) / r146));
		#10; r32 = r221;
		#10; r161 = (((((r79 || 17'h2a79) % $time) !== ($stime + (9'h164 > (r94 * 18'h8a0)))) | (((r104 ^ ((r190 > r53) + $time)) >= r217) > r32)) - r130);
		#10; r10 =  ( & ( ((( ( ! ( r18)) > r102) & ((7'h2c > $time) || (r33 <  ( ! ( ($stime - (((18'h2403 && (((2'h3 <= 7'h46) & r199) + (r138 == ( ( + ( (25'h643f !== 6'h1))) + r82)))) ^ (( ( + (  ( ! ( ((21'h2864 && 4'h9) || (22'h1c12 == 9'he3)))))) || ( ( - ( ((31'h23bf ^ 11'h44f) !== (21'h2257 || 20'h3d63)))) !== (r128 <  ( ! ( (21'h49bf + 25'h936)))))) !== ((($stime ^  ( + ( (7'h52 != 23'h5ce2)))) * ((26'h33f0 | 2'h3) % ( ( ~ ( 24'hafc)) !== r32))) != (r219 == 28'h20f3)))) != r20))))))) | 16'h3a6a)));
		#10; r15 = (24'h31d2 != r30);
		#10; r210 = (r97 | ((8'h4 || r34) ^ (r72 == 11'h724)));
		#10; r214 = ((((( ( ~ ( ( ( & ( 23'h74ba)) > (r92 + (r77 + 4'h1))))) == r26) || ($time != ((12'heb1 <  ( ^ ( ((17'h21be - ($stime >= ((r174 - r230) >= (((30'h1aa7 % 29'h622f) +  ( ! ( 12'h297))) ^ (15'h4020 && r79))))) === r159)))) != $time))) * ((((13'h836 ^ ( ( | ( ((r120 &&  ( + (  ( + ( ((8'he + 30'h2a02) !== r44)))))) % 27'h4d2c))) |  ( & ( (r238 | r214))))) !== (26'h327a != (4'h5 === ( ( ! (  ( & (  ( & ( (((13'h1896 & 22'h33) %  ( + ( 29'h63e4))) + r148))))))) == $time)))) / r173) /  ( - ( r12)))) / r109) && (23'h44f8 > ( ( ! ( $time)) + r205)));
		#10; r182 = ( ( ~ ( 28'h4852)) === 11'h1d2);
		#10; r11 =  ( ^ (  ( ! ( (r142 &&  ( & ( ((r127 <= r51) - 32'h6ebd))))))));
		#10; r221 = 9'h20;
		#10; r97 = ($time + (11'he8 != (( ( ! ( ($time ^ 2'h3))) % (((r175 - (31'h5de9 + 2'h2)) / r70) <= r189)) % ( ( | ( ((r1 || ( ( & ( (5'h11 >= ((7'h3c <= r198) > 16'h5796)))) | 28'h32a)) ^ ((r221 & (($time ^ ((((r220 % (20'h6874 + 4'h0)) !== r219) + 14'h1bd8) / 30'h7574)) + r251)) < (19'h11a4 > r61))))) ===  ( - ( (((r253 + 30'h72b5) < r68) && (((15'h6bf0 > r153) < $stime) !== 6'h20))))))));
		#10; r205 = (((24'h1906 != (( ( ~ (  ( | (  ( - ( $stime)))))) == r74) / 18'h6640)) === r94) + (((27'h1683 == (14'h13fa <  ( & ( r72)))) > r48) * (((((r173 == (4'hd | ((13'ha23 && 1'h1) <=  ( ! ( (9'h1ea ?  ( ~ ( 16'h4ec3)) : ( ( ! (  ( ~ ( (27'h3b76 == 18'h6606))))) * ( ( - ( (23'h3f36 ^ 27'h1521))) % r231)))))))) & ( ( - ( 14'he7b)) <=  ( | (  ( - ( 12'h1d)))))) + r168) <= r217) >= $stime)));
		#10; r231 = (r213 | (((30'h7dd6 && r127) == (r109 | 29'h1794)) != r130));
		#10; r150 =  ( - ( $stime));
		#10; r116 = (r139 > (( ( | ( r219)) <= (29'h25ec &&  ( ! ( 4'h9)))) / ( ( ~ ( r79)) > (r25 ^ 1'h1))));
		#10; r56 = 24'h6d7b;
		#10; r214 =  ( ! (  ( + ( r90))));
		#10; r207 = 19'h5602;
		#10; r116 = ( ( + ( r130)) <= ( ( ^ ( 6'ha)) < r200));
		#10; r220 = (((15'h5ceb + 6'h25) ===  ( ~ ( 11'h1dd))) < r161);
		#10; r10 = r63;
		#10; r63 = $time;
		#10; r214 = r201;
		#10; r225 = $stime;
		#10; r58 = r103;
		#10; r78 = ( ( ! (  ( ! ( r28)))) <= ( ( & (  ( ~ (  ( - ( (r165 && r66))))))) >=  ( ~ ( 6'hd))));
		#10; r243 = 1'h0;
		#10; r25 = ((((21'h9f5 == ((((r24 >= r227) ||  ( ^ ( (r63 ===  ( & ( (r92 >= 21'hc2d))))))) < (32'h71e6 % r124)) - 25'h51f4)) &&  ( ~ ( 5'h17))) != ((r138 || (8'h91 ===  ( & ( (( ( | (  ( | ( r186)))) | r196) !== r186))))) && r103)) + 12'h5cf);
		#10; r175 = (r171 * r99);
		#10; r193 =  ( ~ ( 29'h5007));
		#10; r141 = r64;
		#10; r22 = (5'h11 +  ( - ( ((26'h2b69 ^ $stime) <= (((r129 < (((( ( ! ( 7'h23)) + (4'h5 === (6'h35 >= 24'h20d7))) || (( ( & ( r226)) & (16'h6572 >= (r173 ^ 18'h2888))) - $stime)) ? $stime : 15'hb3d) *  ( ! (  ( | ( r3)))))) < (( ( & ( ((( ( - ( ( ( ~ ( r109)) %  ( ^ (  ( + ( 2'h3))))))) >= ($stime < r136)) ? 7'h5b :  ( & (  ( & ( (((18'h71e * 8'haa) <= (22'h651b - 26'h499e)) | r83)))))) === r134))) == (((20'h65de & (r227 % 7'h63)) >  ( + ( r213))) >= ((9'h18b == 16'h7f14) && ((( ( | ( r78)) < ( ( ~ ( (27'h3ae8 + 31'h566b))) + ($stime >= (16'h55d9 % 17'h7bb4)))) < 28'h3f8b) <= ((r132 != (( ( ^ ( 29'h5761)) ? (6'h5 != 3'h5) : r21) !== r23)) === (2'h0 === r235)))))) == (r49 &&  ( ! ( 9'h11a))))) < r188)))));
		#10; r49 =  ( ^ ( (((((25'h4e96 === r46) && r73) >  ( ^ (  ( | ( ( ( | ( 10'h1b2)) & ((r159 - ( ( & ( r109)) / $time)) >= 14'h1323))))))) - r165) % (r28 > r247))));
		#10; r4 = 30'h3703;
		#10; r165 = r95;
		#10; r39 =  ( + ( (r224 == r178)));
		#10; r248 = $stime;
		#10; r209 = ((12'h657 | ($stime ^  ( ^ ( (r198 != ((22'h1825 + r140) === 26'h5d53)))))) ==  ( ~ ( (( ( & ( ((r21 % (($time | ( ( ! ( (r6 == (((21'h2c09 == 3'h5) == (4'h7 ? 18'h3c25 : 25'h3224)) !== (r13 !== (16'h68df <= 20'haf4)))))) % 9'hc5)) >= $time)) ? 8'hef : (r247 & (r180 ^ ((((16'h31e9 - ($stime & 10'h1bc)) && (18'h7f94 | ($time ? r16 : ((5'hb ? 29'h7896 : 19'h5aba) ^ (19'h52e0 === 1'h0))))) == (((24'h201f !==  ( | (  ( ! ( 5'h1f))))) ||  ( ~ (  ( ~ ( r100))))) / ((r60 ? (r99 || (9'h6 ? 10'h2fe : 27'h72e7)) : (r234 <= (11'h74b % 30'h6ba6))) >  ( & ( ((29'h4113 !== 29'h4226) && (5'h1e > 15'h3bb0))))))) != ( ( + ( ((1'h1 - 1'h1) >= (r31 * ($time ? 22'h7283 : (10'h25c == 1'h0)))))) & (r57 === (9'h1e9 < r56))))))))) >= 7'h17) != r163))));
		#10; r1 = (r78 % r79);
		#10; r101 = ( ( ! ( (((r143 - 30'h78e0) / (14'h1c2e - (((( ( ~ ( 27'h5102)) !== 23'h5656) *  ( + ( (r127 >= (((((31'h4150 == 9'h7f) ? (21'h40b0 >= 1'h1) : 20'h7e04) >=  ( | ( 31'h6fed))) ? ( ( + ( r11)) && (15'h1543 && (8'h45 < 24'h382b))) : r189) > (r201 <= r171)))))) && ($stime > r42)) &&  ( & ( 14'h39ec))))) == r110))) === ((($time /  ( - (  ( ! (  ( + ( 1'h1))))))) & r199) !== 12'h112));
		#10; r111 = $time;
		#10; r58 = r34;
		#10; r1 = (21'h4628 & (r206 >= r167));
		#10; r130 = (( ( ^ ( r212)) + r148) !== ((r51 !==  ( + (  ( ~ ( ((8'h68 == $stime) >  ( & ( $time)))))))) || 6'h0));
		#10; r12 = (( ( & ( ( ( - ( (((r233 && (r155 || r64)) > (r224 != ((19'h1e80 * (24'h7122 & ( ( ! ( r79)) | (r81 >= r68)))) != 11'h3de))) ? ((r139 > (21'h58b4 < (($time - ($time | 1'h0)) === (((14'hf05 | 9'h90) ? (r180 -  ( - (  ( ~ ( 4'h3))))) :  ( - ( 12'h8e9))) >= ((9'h195 > ((13'h19a8 < 23'h5a73) && 7'h21)) && $stime))))) ^ r46) : ((r171 !== ((((9'h120 != (2'h0 %  ( + ( r237)))) &  ( ! ( 3'h6))) || (( ( & ( (31'h7 || 23'h777a))) !==  ( - ( (r102 + (1'h0 + 26'h4b6a))))) & $time)) * r78)) !==  ( ^ ( $stime)))))) != 13'haee))) ? r59 : (29'h3976 / r181)) % r221);
		#10; r246 = r187;
		#10; r122 = 32'h7516;
		#10; r63 = r192;
		#10; r68 = 21'h5966;
		#10; r221 = (( ( - ( (r154 === 2'h3))) && ( ( ~ (  ( - ( $stime)))) > $stime)) ^ ((27'h464f <= r132) < 24'h4012));
		#10; r179 = r107;
		#10; r15 = 26'h1958;
		#10; r27 = (r197 != r242);
		#10; r251 = (2'h1 <= 7'h69);
		#10; r252 = (r50 <= r231);
		#10; r228 = r192;
		#10; r181 = r218;
		#10; r129 = ((r187 & (($time || (r85 >  ( ~ ( r13)))) > 32'h2b02)) | ($stime !== ( ( ^ ( r164)) +  ( ^ (  ( & ( ((((((( ( - ( 9'h133)) - r240) && 10'h1e0) <= 12'h481) >= ( ( ~ ( (r78 !== (r132 | r63)))) %  ( + (  ( - ( ((r159 &  ( & ( 29'h376e))) >= ((1'h1 || 30'h4e92) && (19'h1691 & 26'h2629))))))))) * (r200 == ((r202 > (((r83 % (14'h2086 == 12'h1ca)) >  ( & ( r246))) <= (((6'h7 + 23'h27fb) ? (1'h0 !== 15'h3dbc) : $time) - (r117 <= (9'hcb != 19'h31ef))))) ? 2'h0 : ( ( - ( 8'hb7)) || r65)))) ? ((r92 != ( ( - ( ( ( ! ( 25'hc76)) && 17'h27e3))) >= ($time == (r196 ? (((19'h842 != 17'h44a4) &&  ( ^ ( 3'h3))) / r124) : 1'h1)))) *  ( ^ ( r17))) : (10'h300 <= (($time | (r161 !== $time)) - r55))) &  ( + (  ( + ( $time))))))))))));
		#10; r69 = (( ( ! ( r209)) != 27'h73e0) / 30'h5ff5);
		#10; r36 =  ( ^ ( (($stime % 22'h7f73) /  ( ! ( (r60 / r187))))));
		#10; r195 = r61;
		#10; r148 =  ( ! ( ((r1 != r174) & r111)));
		#10; r61 = r232;
		#10; r86 = (11'h627 / (( ( | ( r110)) <  ( ^ ( 25'he53))) > (((( ( & ( (20'h1ed3 - 4'h9))) <  ( ^ (  ( & ( 15'h48a3))))) | ((r73 % r163) && (((($stime !== ((r195 || ((18'h61d8 | (2'h2 + 32'h6491)) ? ((9'h1bd & 21'hdab) * (16'h597b == 5'h15)) : 27'h1e00)) & r87)) ? ((16'h6477 | r71) > ( ( ! ( 17'h49a5)) == r179)) : (( ( - ( ( ( ! (  ( & ( 26'h2396)))) + (19'h3d37 & (30'h1edf === 18'h2788))))) && (((r165 != 14'h13b0) ? r203 : $time) >= (r242 + r68))) <= r147)) ?  ( ~ ( $time)) : (r189 + r151)) >= 8'h98))) === 25'h4203) ? $time : ((29'h133a ^  ( - ( (r137 !== 6'h1d)))) || ((( ( + ( r50)) || ((r216 === 32'h7fe7) >= (9'h13d >= r229))) &&  ( + ( 19'h2336))) & r246)))));
		#10; r19 = (r85 | (24'h5e3d ^  ( ^ ( (r246 == (18'h6068 &  ( & ( r152))))))));
		#10; r4 =  ( + ( $time));
		#10; r152 = ((( ( - ( r140)) | ((1'h0 ? (1'h1 && r199) : (( ( + ( r212)) == r72) * ((r4 !== 5'h3) > (($stime >= 31'h742c) <= (13'h131c < r213))))) > (r246 || ((r116 < (((r189 <  ( & ( ($stime === ( ( ^ ( r100)) | r189))))) !== ((r96 | ( ( ^ ( (r40 & r20))) * r167)) - (((r219 || 5'ha) === r185) != 20'h34fd))) | 17'h2d95)) + (( ( + ( (r114 % 25'hab5))) <= (( ( | ( r206)) ||  ( & ( ((18'h2670 &  ( + (  ( & ( 14'h24d9))))) ? (14'h3df < (r253 | 19'h514e)) : (r5 * ((29'h88e != 15'h202c) <= (25'h7dd4 || 21'h4915))))))) === 7'h7d)) === 32'h2450))))) / r139) >=  ( ^ ( ( ( ^ (  ( | ( 31'hc9a)))) >= 27'h5ce1))));
		#10; r83 = r149;
		#10; r106 = (((r142 + (18'hff6 - r189)) ?  ( & ( (r109 && 30'hb4f))) :  ( - (  ( | (  ( | ( r115))))))) <= r180);
		#10; r227 =  ( ! (  ( ! ( ($stime / ((r194 * 26'h6311) === ((r105 % r76) != ((r79 != (1'h0 || (((2'h3 >=  ( ^ ( 4'h4))) - 23'h5b50) > r48))) ^ 27'h702))))))));
		#10; r38 = r32;
		#10; r177 = (r151 ^  ( & ( r53)));
		#10; r132 = r245;
		#10; r135 =  ( + ( (r141 - ((r169 != r178) !==  ( | ( (r241 !=  ( & ( ((r102 &  ( ~ (  ( ! ( r18))))) ^ r25))))))))));
		#10; r121 =  ( | ( 18'h61eb));
		#10; r253 = (((r123 >= 13'h18f9) & 26'h1e42) ===  ( + ( (r185 < r245))));
		#10; r58 = r52;
		#10; r1 = (( ( - ( 21'h3df1)) === r43) && r195);
		#10; r180 = ( ( | (  ( + ( 23'h51f6)))) | $time);
		#10; r147 = r50;
		#10; r212 = (r48 /  ( | ( ( ( - (  ( & ( (r78 & r199))))) ^ (((r190 !=  ( & ( (r11 * (( ( - ( (($stime <= ((5'hd ? 11'h55e : 21'h7496) === (6'h23 % 15'h406b))) || r52))) / $time) > 18'h68f1))))) - ((($stime == r49) & r191) > (( ( ^ ( (13'h11e6 - 2'h0))) === (((8'h77 > ((( ( & ( 18'h6c31)) + r247) + (r154 <  ( ! ( 15'h2dda)))) >= ( ( - ( $time)) ^ ((4'h0 * 19'h3e9c) | r11)))) != (r70 != ((((18'h2d84 != 2'h3) != r202) / ((29'hf27 !== 29'h5512) + r43)) !== (18'h1db <  ( & ( r221)))))) / r255)) ||  ( + ( (r32 + (r106 - r168))))))) || $time)))));
		#10; r140 = (r210 - ((((r91 >= 25'h6118) & r15) >= $time) - (((((23'h4c9c ? r228 : ( ( + ( 27'h4433)) == (r117 == ((($stime | (($stime |  ( & ( 23'h52a9))) === (r138 || r157))) === r106) * (r190 != $stime))))) |  ( + ( r200))) - 28'h7a48) === 12'h1be) / ((r45 - ($stime + 4'h2)) != (( ( + ( (27'h7bf7 | (((27'h1e92 % 5'h17) ? 17'h4f68 : r240) >=  ( + ( ( ( & (  ( - ( ((27'h6ca1 | 4'h5) ? (1'h0 ? 15'h551a : 19'h3554) : (2'h1 ^ 24'h62bd)))))) >  ( ~ ( r248))))))))) ^ r123) * r183)))));
		#10; r116 = ((($time * (7'hd !== $stime)) >= 12'h528) + 2'h2);
		#10; r16 = r182;
		#10; r188 =  ( - ( 15'haa4));
		#10; r235 = ($stime ?  ( ~ ( (30'h4340 > $stime))) : r134);
		#10; r206 = (21'h355e && 16'h3c42);
		#10; r32 =  ( - ( (22'h3162 < ((r236 === 17'h4e9f) !=  ( ~ ( r231))))));
		#10; r2 = 4'h4;
		#10; r227 =  ( - (  ( ~ ( r70))));
		#10; r123 = r227;
		#10; r52 = 11'h62c;
		#10; r187 =  ( & ( (28'h554a !== r129)));
		#10; r15 =  ( ! (  ( - ( ((14'h23b | ((24'h5d96 < ( ( ^ ( r81)) % ((26'h13a2 - (((10'h2d4 <= (((7'h1d < 23'h784b) <= 2'h0) <= r41)) % ( ( - ( r76)) >= (7'h54 || ((20'h667a * 7'h4a) != (16'h3c25 | 18'h732))))) ? (r125 ? ( ( ^ ( (r6 == (32'h1414 + 30'h61ef)))) & (r75 != 27'h17c1)) : (r157 - ($stime / ( ( ^ ( 1'h1)) ?  ( ! ( 22'h5660)) : r112)))) : (r244 & ((1'h0 >= r112) === ((r203 >= r3) + ( ( | ( 12'h2a8)) < (30'h838 + 17'hb72))))))) - r84))) | ( ( ^ ( ((23'h151 / ( ( ~ ( ( ( ^ ( ((6'h29 - 11'h624) % $stime))) +  ( ! ( ((32'h5711 ? 3'h6 : 28'h4941) % (19'haad === 12'h299))))))) + 14'h340c)) ^ 12'he4f))) !== r64))) | (( ( | ( ( ( ! ( ( ( & ( ( ( | (  ( | ( 9'h1a2)))) /  ( ^ ( (11'h15b ? (r141 == $time) :  ( | ( r242)))))))) == (24'h338 == r170)))) !== 20'h28f8))) <= (((r75 >=  ( ~ ( ((( ( & ( 16'h5800)) &&  ( ~ ( r186))) & ((r215 / r60) <= (((32'h1ce6 | 15'h3e47) <= (1'h0 <= 29'h3f9c)) !== ((23'h5d5d <= 23'ha77) | (9'h20 < 22'h43a4))))) % ((9'h39 + r179) || r82))))) -  ( ~ ( r243))) > $stime)) ? ((r105 > (r217 + 27'h2e68)) ? r223 : r81) : r31))))));
		#10; r228 = r194;
		#10; r187 = 7'h29;
		#10; r109 = ( ( ^ ( ((13'h1f6 >= r210) + r112))) > r235);
		#10; r121 = 13'h5bb;
		#10; r213 = ((r30 * 18'h2845) ===  ( ! ( r237)));
		#10; r180 = ((r241 | (((r106 - (( ( + (  ( ~ (  ( + ( 28'he39)))))) !==  ( - ( (($stime | ($stime != (((r139 % r97) !== r94) >= r251))) ^ r45)))) | r97)) === (r79 < ((r109 * 2'h0) !==  ( & ( 27'h3293))))) / (((r238 + 15'h60cb) == ((( ( + (  ( | ( r65)))) <=  ( & ( 29'h7fa4))) > (($stime | (((r24 <  ( - ( 10'h116))) % ((($stime >= (14'h2dac | 4'h2)) / (5'h1 && (11'h68e != 12'hfd))) | r57)) - r252)) ? 30'h2533 : r239)) < r117)) === r175))) % 25'h5022);
		#10; r7 = (( ( | ( (15'h7910 &&  ( & ( (r66 <= r105)))))) < (29'h6770 %  ( ^ ( r24)))) + (r27 - (($time * (( ( ~ ( ( ( & ( r72)) ||  ( ~ ( ((16'h613e ? (6'h18 + r105) : ((r58 ^ ( ( - ( 1'h0)) > (15'hd9d | 12'h8d8))) > ($time === r11))) + ((r60 + r170) >= (30'h109b ^  ( - (  ( + ( (19'h3346 ? 12'hf5 : 21'h2119))))))))))))) < 5'hf) - $time)) !==  ( ~ ( ((r246 >= (((r90 - 14'h34ad) !=  ( | ( 25'h6134))) && ( ( ! ( ( ( | (  ( | ( (r152 | r232))))) |  ( ~ ( (r196 || r35)))))) ||  ( - (  ( & ( ((r73 >=  ( & ( $time))) ||  ( - ( (23'h1d25 !==  ( + ( (20'h672d === 24'h194b)))))))))))))) == ( ( & ( r34)) !== (r30 /  ( & ( (( ( ^ ( 17'h6d41)) ?  ( + (  ( ~ ( (11'h77f || ((1'h0 - 31'h185d) == (28'h1b96 ^ 15'h2a2a))))))) : $stime) != ((19'h7835 ==  ( ! ( 32'h4eb6))) ||  ( ! ( (( ( ^ ( $time)) ^  ( + ( (16'h1f16 + 22'h17f)))) == r118)))))))))))))));
		#10; r21 = 24'h1fe8;
		#10; r145 = (( ( - ( 17'h64a4)) !== ((r131 > (r109 | ( ( ~ ( 14'hd50)) + (r228 !== (( ( ~ ( ((29'hc3f - (( ( | ( 27'h6286)) <= 18'h6b93) === 31'h2432)) && ($stime || ( ( | ( 23'h35a)) <= 32'h496))))) && r113) == r175))))) <= r252)) && r171);
		#10; r210 =  ( - ( (r171 != (r235 > r32))));
		#10; r212 =  ( & (  ( ~ ( ((r90 != r45) & 11'h491)))));
		#10; r158 =  ( - ( 14'h3cb));
		#10; r152 = (r137 ==  ( & (  ( + (  ( ~ ( 18'h3802)))))));
		#10; r152 = r114;
		#10; r28 = (r72 % r210);
		#10; r69 =  ( & ( ( ( - (  ( ~ ( (( ( ^ ( (((((22'h7b4e < ( ( & ( (7'hb > 31'h50d8))) ^ (4'hb / (17'h3b5d == 7'hf)))) & r220) % (8'h4e <  ( ! ( 18'h2d17)))) - r130) * (16'h4fd5 * ((( ( ^ ( 24'h716d)) &&  ( ! ( r221))) >= $stime) == (31'h4a6f > ((r24 & ( ( ^ ( 30'h309)) <= (29'h475 == 28'h2d97))) >=  ( & ( ((30'h151f <= 22'h6762) * 17'h646b)))))))))) - ( ( | ( r45)) * r211)) == ((r114 / $stime) === (21'h2915 !=  ( ~ (  ( ! ( $time))))))))))) == ((r197 || 27'h73e0) <= 14'h3d7))));
		#10; r60 = (( ( | ( r187)) == ( ( - ( r55)) + (((11'h335 > (r232 != r5)) == (r89 ? ( ( | ( $time)) !== r6) : ((22'h6cc5 && (9'h161 <= $stime)) <= $stime))) <= r123))) / (((( ( ~ ( $stime)) >=  ( | ( r221))) <  ( - ( r115))) !== ( ( ! ( (( ( ^ ( (( ( & ( r95)) + (13'h49d <  ( | ( 18'h1a82)))) !== ((r78 != (r34 >= ( ( ! ( (14'h588 | 16'h507))) && (1'h1 > 12'hbfd)))) && (r91 + r249))))) !==  ( ^ ( ( ( | ( r205)) == r71)))) == 15'h113d))) === 32'h60ad)) /  ( + (  ( - ( 15'h7b84))))));
		#10; r213 = ( ( + ( 3'h0)) / (8'hc6 < r26));
		#10; r27 = 19'h54d6;
		#10; r235 = (10'h2ce || (14'h18b5 * ((($stime & ( ( ~ (  ( ^ ( (((((r39 ? ($stime % 7'h68) : ( ( ^ ( 7'h38)) || (14'h99b % 24'h613f))) != (r116 < r163)) | r154) ?  ( - ( 22'h2d1e)) : 12'hf49) - ((((((19'hee0 + 25'h4274) === r189) + 21'h1c66) * 25'h2b72) &&  ( ~ ( (( ( ~ ( 18'h4339)) & 6'h3e) %  ( + ( (10'h218 | 19'h4ea1))))))) == ( ( - ( r117)) | ( ( | ( r118)) | (r63 !==  ( + (  ( ~ ( 27'h3763))))))))))))) < r82)) & r142) ==  ( + ( (23'h74ab &&  ( ~ ( r108))))))));
		#10; r3 = 24'h3a7b;
		#10; r60 = ( ( ! ( 22'h5ca)) |  ( ! ( (r38 / (r0 ^ ((30'h7151 ^ ( ( + ( 1'h0)) ^ (4'hc || (r49 > (14'h1287 %  ( | ( (3'h2 !== (((26'h1516 != 4'ha) + 19'h7343) < (r225 *  ( & ( 27'h380d)))))))))))) < r55))))));
		#10; r209 = $stime;
		#10; r88 = 30'h47b0;
		#10; r190 = ( ( - ( r25)) != (r230 % r145));
		#10; r242 = (((r31 ^ r98) ^ (( ( | ( r110)) < ((( ( - ( ((( ( | ( (r147 != r193))) | 15'h2197) &&  ( ~ ( ((((9'h1b / 3'h6) - (16'h66b5 !== 13'h15aa)) <= (r188 || (24'h1e3f >= 30'h41da))) <= (r181 / ((11'h317 - 30'h7563) <= (32'h1a3a && 8'h20))))))) * $stime))) ?  ( & (  ( & ( 21'h5bc5)))) : (3'h2 - 10'h332)) % r29) <= r182)) == r131)) ^ (24'h3d27 && (28'h3b13 !== 20'h1322)));
		#10; r227 = 23'h11c3;
		#10; r242 = ((21'h5910 == (19'h6d6f -  ( ! (  ( | ( r100)))))) <=  ( + ( (r208 - ( ( ^ (  ( & (  ( ~ ( r170)))))) / (((r216 && r115) != (r68 ? (1'h1 * r149) : 2'h3)) && r233))))));
		#10; r178 = r186;
		#10; r44 = ( ( - ( r213)) && ((r59 % r72) / r65));
		#10; r26 =  ( - ( r97));
		#10; r120 = $time;
		#10; r251 = r73;
		#10; r78 = 25'h4661;
		#10; r105 = ((27'h3d8e | r115) || 19'h65b7);
		#10; r212 = (11'h727 > r67);
		#10; r198 = r128;
		#10; r59 =  ( + ( r140));
		#10; r125 = 19'h6ff4;
		#10; r99 = ( ( + ( r41)) === 30'h295e);
		#10; r197 = r17;
		#10; r5 = (r172 === r139);
		#10; r252 = (((17'h64d7 ^ 4'hd) + ( ( | ( ((13'h19cb && r127) %  ( + ( (25'h69d4 >=  ( + ( 17'h956)))))))) > (((( ( ~ ( 18'h5835)) | ((((r63 | 22'h33eb) < 19'h7c40) | 22'h1c7e) % ( ( - ( (r77 >= ($stime ? 21'h1762 : (((4'ha > 14'h2fb0) < 16'h2d72) |  ( - (  ( ! ( 32'h2f02))))))))) +  ( + ( ( ( ~ ( (r60 ? $time : r244))) >= 28'h67c5)))))) <= (r106 & 32'h28a6)) != r242) / 6'h39))) ==  ( & ( 9'h1e2)));
		#10; r58 = r119;
		#10; r102 = 17'h597e;
		#10; r148 = r206;
		#10; r22 = (r194 ^  ( | ( 26'h249c)));
		#10; r133 = (((r34 | (20'h12d2 === r166)) != ($stime !==  ( ^ ( (($time == r53) ==  ( - ( 4'h6))))))) !==  ( ~ ( 5'h13)));
		#10; r182 = r102;
		#10; r165 = ((r60 / r30) % r33);
		#10; r20 = ( ( + ( r17)) != r90);
		#10; r102 = (((r105 - (20'h3e12 < 24'h5669)) > (((21'h12ed != ( ( | ( (r82 > ( ( ! (  ( & ( (r187 <  ( + ( ((12'haa1 === 4'h8) + (32'h2954 % 11'h3be))))))))) + (21'h74de * 3'h4))))) -  ( ~ ( 16'h6332)))) / ((r178 ||  ( - ( 30'h6f10))) | 31'h5072)) ? ( ( ~ ( (( ( ~ ( (r197 >= $time))) >= r254) > (r51 ^ 5'h5)))) !== ((((r82 > ((r40 != (r68 < ((((23'ha77 * 20'h39dc) * (31'h87c / 16'h5e84)) | (32'h666b % (13'haac >= 31'h757c))) === 6'h5))) || (r254 <= ((((7'h3c / r179) + r196) != r61) !== ((11'h27e - r0) <= (($stime >= r0) / 15'h2676)))))) !== r49) *  ( - ( ((r106 &&  ( ~ ( 23'h50ed))) >= (11'h77e <  ( ^ (  ( ~ ( 2'h1))))))))) !== $time)) : ((r242 >= ($time !== (r169 > (18'h129 == 32'h4fe8)))) <  ( & ( (((32'h925 || r56) ? r180 : 18'h5ecc) === (( ( - ( 14'h23fa)) & (r203 ==  ( | ( (17'h78cf <=  ( - ( (r223 | ((1'h1 < 14'h251f) ? 5'h1c : (28'h52ce >= 27'h1c52)))))))))) - r233))))))) <= (( ( ~ (  ( ^ ( ($stime / r49))))) + r27) !== $time));
		#10; r21 = ((r8 ? 2'h1 : (( ( ~ ( (r82 + $time))) < r44) | r98)) / r188);
		#10; r4 = r126;
		#10; r91 = 11'h2c3;
		#10; r113 = 18'h3ed2;
		#10; r47 = r29;
		#10; r128 = ( ( | ( 9'h35)) ^ 27'h35ad);
		#10; r120 = r110;
		#10; r54 = ((r68 !==  ( ! ( r28))) == (25'h571a & ( ( - ( ((r161 & 23'h6f59) !== ((r150 || 18'h6a2f) | 5'h19)))) ||  ( ~ (  ( ~ ( ( ( ~ ( $stime)) ^ r68))))))));
		#10; r246 = ((23'h18f0 ^ r230) + ((((18'h4781 ^ r148) > (((r247 - 2'h3) == $stime) >= ((((r170 || (r209 !== ((6'h18 % r248) === r170))) > r2) || ((((4'h5 + ((( ( + ( 4'h9)) & (31'h206f <= 32'h74e0)) <= ($time / (12'ha4e !== 12'h1b8))) > $stime)) === ($time > (((r98 <= r156) | r171) ||  ( - ( ((2'h0 > 29'h52a5) - r155)))))) & (r80 ^ $stime)) == r118)) == ((r122 % ( ( ^ ( 9'h61)) ===  ( ^ (  ( & ( r57)))))) ^ ((((r168 || ((r149 > (r65 -  ( | ( 16'h3096)))) >= $stime)) <  ( | ( (20'h30d5 - r250)))) != (((( ( | ( 8'h72)) ^ r193) <  ( & ( (17'h13cf ^ (18'h57e0 <= 5'h1d))))) * r163) * (9'h1ff === ($time | 29'h1f07)))) > ($stime ||  ( | (  ( ^ ( ($stime > (r182 >= $time)))))))))))) === ((32'h7235 +  ( + ( r63))) != (25'h5617 !== r193))) > (26'h3b84 <= r37)));
		#10; r61 = ((( ( + (  ( - (  ( | ( (9'h123 < ((((r131 == $stime) !== r221) ^ $time) >= (26'h7d2b && (16'h4c88 === 28'h630e)))))))))) / (29'h2ad5 <=  ( + ( ((r198 * ((r25 * (r33 + 4'h9)) <= r172)) != ((r173 >= 27'h16a3) < (r24 != 10'h27d))))))) & ($time / ($stime &&  ( + ( (23'h2212 ? (r86 <=  ( ^ ( (10'h2f2 > (r126 / 30'hc28))))) : (r16 |  ( - (  ( + ( (r0 <= (((14'h3e2f <= r129) < r115) !==  ( - ( r156))))))))))))))) || 20'h118);
		#10; r132 =  ( ^ ( r44));
		#10; r100 = (r14 ==  ( | ( ((r236 != r163) & $stime))));
		#10; r46 = (30'hc90 - r136);
		#10; r99 = (r38 + (r75 &&  ( ^ ( 1'h1))));
		#10; r110 = ((5'h1c + 12'hd0d) ? (( ( ! ( r29)) |  ( ~ ( (5'h4 < (8'h1a != 9'h11))))) == r103) :  ( & ( ((((r69 &  ( & (  ( & ( r222))))) % ((6'h39 <  ( + ( 10'hd3))) === r11)) ? (r252 === 6'h25) :  ( ^ ( (( ( ! ( 20'h774a)) | 30'h2641) |  ( | ( (((5'h4 !== r29) == ((r204 ^ r33) || 14'h465)) > (r161 <= r169)))))))) >= r231))));
		#10; r227 = (r186 ^ (($stime /  ( - ( ((((30'h5a52 != (( ( ! ( 8'h49)) === (r202 | 8'h31)) == r148)) <=  ( - ( (11'h388 & 11'h6fb)))) === r104) < r226)))) + 1'h1));
		#10; r62 = 19'h4ab;
		#10; r231 = r234;
		#10; r111 = (r230 * $time);
		#10; r25 = $time;
		#10; r186 = ( ( ! (  ( | ( $time)))) ^ r243);
		#10; r235 = r235;
		#10; r38 =  ( & ( (( ( ! (  ( ! ( 15'h298c)))) / (((r103 % (5'ha >= r102)) ^ 16'h6162) / 24'h2416)) < ( ( - ( r135)) &&  ( & ( r148))))));
		#10; r49 = ((( ( ~ ( $time)) < (r116 % 23'h2cb1)) > (20'h4454 ?  ( | ( (21'h198e | $stime))) : r116)) ^ (r55 ? r252 :  ( ! ( (r154 ?  ( ^ ( 16'h6adc)) : (23'h284 > (( ( - (  ( - ( 27'h2f79)))) <= r130) <= (( ( | (  ( ~ ( $stime)))) !== ((r25 ^ r1) === r199)) !== ($stime > ( ( & ( 23'h2b4)) < (r247 || 10'h190)))))))))));
		#10; r169 = (((r12 | r195) > $stime) * ( ( + (  ( - ( (r20 >= (13'h508 === 18'h11fc)))))) ||  ( ! ( 18'h2923))));
		#10; r199 = $time;
		#10; r224 =  ( ~ ( ((23'h4d5 & r216) && r228)));
		#10; r46 = 23'h79a5;
		#10; r94 = 6'h1e;
		#10; r46 = r181;
		#10; r103 = (( ( ~ ( (((8'he6 - r129) < ((r204 + (10'h139 % r112)) < r75)) | ((r96 >= 25'h4652) != (r216 * r46))))) >  ( ! ( ((20'h7cc1 < 19'h1460) || r74)))) & r190);
		#10; r61 = ( ( & ( (r33 < (r53 <= r38)))) !== r135);
		#10; r12 =  ( + ( (( ( ! ( $stime)) || 3'h7) + (( ( ~ ( (3'h4 + ((r189 ? (30'hc61 >  ( - ( (7'h21 ? ((((29'h5467 | 3'h2) || (31'h2f57 >= 11'h760)) ^ ((4'h0 & 16'h5c22) * 7'h39)) ===  ( + ( $time))) : (21'h546f > (1'h1 | ( ( - ( 4'h5)) *  ( - ( 26'h144))))))))) :  ( ! ( r186))) === r251)))) + r49) | r241))));
		#10; r173 =  ( - ( r247));
		#10; r65 = $time;
		#10; r57 = 10'h120;
		#10; r230 = ( ( ~ ( (r203 * r115))) ? r16 :  ( ~ (  ( ^ ( r204)))));
		#10; r201 = (r58 <= r7);
		#10; r63 = r217;
		#10; r93 = (17'h70ab - ( ( ~ ( 5'hd)) ^ (( ( ~ ( ((( ( & ( ((17'h63e4 % ((((19'h70fc * 10'h1fa) === 23'h5ba5) - 25'h830) ^ r254)) - 1'h0))) !=  ( ^ ( (((( ( - ( r27)) & r177) % r226) / 8'h24) * r209)))) | 30'h1439) != 22'h7b4b))) / (r51 + r174)) <=  ( + ( r65)))));
		#10; r243 = 8'heb;
		#10; r97 = ( ( & ( ((r126 % 15'h4856) <  ( + ( r14))))) !== r25);
		#10; r233 = 18'h5ffb;
		#10; r157 = (r172 >= 29'h2fdf);
		#10; r22 =  ( | ( 5'hd));
		#10; r231 = r89;
		#10; r144 = 26'hd4f;
		#10; r83 = $stime;
		#10; r108 = 12'hbe2;
		#10; r45 = (r215 === (( ( + ( 30'h2e06)) <= r205) == (( ( | ( r142)) !== 13'h1108) == ( ( - (  ( ^ ( r253)))) == 31'h19c2))));
		#10; r22 = r84;
		#10; r251 = ((( ( & (  ( ! ( r75)))) <= r183) * r79) < ((1'h0 !== 29'h11fc) !== r124));
		#10; r216 = (r168 &&  ( + ( r70)));
		#10; r104 = (28'h322b ? $time : (r71 - ((r27 ? ( ( ! ( 18'h42a9)) < ($time === (12'hfca * (13'haae <= ( ( + (  ( - ( r86)))) + ( ( ^ ( 3'h3)) == r20)))))) : r86) | ((((22'h689 + ((11'h164 ? r93 : (31'h5fb0 /  ( ~ ( ((((13'h228 === 30'h1aac) && (32'h6fa6 / 13'hce9)) - ((2'h0 & 14'h32e3) < (5'h5 > 9'h1f4))) && 14'h2bcb))))) % (17'h2ebf ? 2'h3 :  ( & ( r237))))) <= ((r84 * ( ( | ( r121)) || r158)) * r54)) /  ( ! ( r74))) != r209))));
		#10; r195 = (r229 ^ (r139 - ( ( ! (  ( - ( r80)))) !== ((10'h17b >= (r243 > (r164 != 2'h1))) < 5'hd))));
		#10; r234 = (r252 ^ (((r76 | r123) / r202) && r219));
		#10; r235 =  ( | ( r121));
		#10; r163 = ( ( ! ( $time)) != (2'h3 ? r30 : (r38 % 26'h781f)));
		#10; r118 =  ( & ( r48));
		#10; r27 =  ( | (  ( ! ( r110))));
		#10; r226 = (r163 * 20'h3fca);
		#10; r170 = (r217 && r180);
		#10; r22 = ((r234 > 27'h2e9d) / 6'h35);
		#10; r158 = (1'h1 === 9'h122);
		#10; r83 = r244;
		#10; r189 = r11;
		#10; r233 =  ( & ( (4'h6 <= (((r254 / r74) + (r104 < ((31'h6871 !== ( ( ^ ( (r235 === $time))) ? (($time % r158) && (23'h4695 >  ( ~ ( 9'h165)))) : r225)) || (( ( + ( r138)) - r213) < (r43 ^  ( | ( r91))))))) >= ($time + (r186 ? 27'h3860 : r182))))));
		#10; r29 = (((((5'hf + (r171 == $stime)) !== (30'h4076 === (((11'h1e2 <= (17'h234d ||  ( | ( 20'h6b6b)))) < r173) || 24'h400b))) | r90) % (22'h620b <= ((5'h4 * 19'h67f7) > r168))) &  ( + ( $stime)));
		#10; r251 = r250;
		#10; r192 = r214;
		#10; r126 = r114;
		#10; r91 = (25'h4e2b + ((((r213 ||  ( ! ( (r79 % r144)))) !== (r251 ^ r127)) % 5'h1) == ( ( ^ ( 7'h2e)) * r254)));
		#10; r156 = 23'h3c0;
		#10; r224 = r158;
		#10; r255 = (( ( ! (  ( & (  ( | ( r88)))))) == r179) >= (r137 || 31'h4d5f));
		#10; r69 = (((r77 || 15'h4f09) ^ ((( ( ~ ( ((r190 ? 4'h6 : ((r135 && ((r151 || 13'hb64) -  ( ! ( (r38 % r115))))) != r54)) | ((((r8 + ( ( ~ ( ((22'h50de >= 4'h5) || (10'h3af !== 10'h188)))) < (((13'h8ac * 28'h65db) ^  ( - ( 32'h108))) - ((14'h13c7 == 28'h60f6) !== r253)))) < ($time - ((r11 &  ( - ( (17'h29f6 == 25'h56c9)))) == (5'hb > r51)))) <= r88) < 15'h7b0f)))) *  ( - ( r197))) & ( ( - ( r234)) >= ((((12'h529 < ((20'h486a <= (8'hbb == (r4 !== r114))) > ((r68 == 1'h0) - ((r172 ^ r108) >= ( ( ~ ( (22'h5e34 + 25'h35ec))) == r26))))) ? (r30 *  ( ! ( (r65 != (((r105 | 3'h3) - ((3'h5 - 10'h315) - 25'h4df9)) | ((9'h1e6 ^ 21'h2aa2) - ((13'h17bb >= 21'h7f98) == $time))))))) : 17'h7c99) / ((r174 | ((r61 != (r233 ==  ( + ( ( ( | ( 20'h6357)) !== r173))))) != r219)) % (24'h6372 ===  ( | ( (((((15'h5a99 / 19'h2862) || (4'h0 & 28'h5982)) == r65) && $time) / (( ( + ( (12'h15f + 8'h97))) < r96) != (r100 <= (r142 >= 3'h3))))))))) * (( ( - ( (r30 !==  ( | ( ((((2'h0 | 9'h61) && (14'h3841 && 11'h620)) !== (r236 / r38)) && r68)))))) & r95) ^  ( ~ ( r92)))))) <  ( + ( (r76 === $stime))))) ==  ( ! (  ( ^ ( (((31'h5d2f >= r92) - (($stime >= r103) < ((r128 | 23'h22f1) % (20'h47b3 < ($time ===  ( | ( r180))))))) / 25'hb6e))))));
		#10; r233 = ((r44 >=  ( ! (  ( & ( (21'h38fd || (r106 % (r184 &  ( ~ ( (r158 & r174))))))))))) / (7'h38 % (r100 & ((r11 - r201) ? (r130 +  ( ^ ( $stime))) : (( ( ~ ( (1'h1 ^ r76))) -  ( & ( (3'h0 >= ( ( & ( r50)) != ($stime | r49)))))) + (30'h6282 * 29'hfe6))))));
		#10; r214 = (30'h1532 / ((((r137 && (r27 - $time)) | ((r222 >= ((r101 ?  ( & ( (( ( + ( r93)) &  ( ~ (  ( ~ ( ((12'ha8d && 10'h1b2) > r62)))))) +  ( ~ ( r201))))) : r235) !== (($stime ^  ( | ( r92))) & (20'h3e39 > ((32'h39ff - (r181 === r17)) || r160))))) ^ (32'h4120 *  ( - ( (22'h7d08 < ((32'h74fd != (( ( - ( 4'he)) >= ((23'h7cee <= r20) &  ( + ( (20'h4711 / 32'h1bb6))))) + ((((21'h2fec === 13'hd08) === 7'h22) <= ( ( ! ( 17'h6a6)) == r109)) | ((9'h1c + (1'h0 | 29'h4e54)) >= $time)))) - 29'h5ff4))))))) !== r237) / 10'h256));
		#10; r26 = (27'h3abb & ($stime * r112));
		#10; r28 = (r212 < 4'hd);
		#10; r128 = r109;
		#10; r59 = $time;
		#10; r180 = r37;
		#10; r109 = 6'h10;
		#10; r80 = (r0 > r215);
		#10; r26 = 2'h1;
		#10; r185 = (7'h76 !== ((((r221 - (((r159 !==  ( ~ ( 16'h110b))) || (r133 % $stime)) & (r66 - 30'h5f20))) !== 8'h99) - r170) == (25'h345f !== (r78 ^ ( ( + (  ( ^ (  ( - ( (r196 ^ $time))))))) !== (5'h1 && (10'hee - (19'h4256 ^ r246))))))));
		#10; r146 = 26'h1c07;
		#10; r69 =  ( + ( r129));
		#10; r187 = (((r245 |  ( & ( 6'h32))) == 28'h34e2) || r128);
		#10; r38 = $stime;
		#10; r233 =  ( ^ ( 18'h57d6));
		#10; r174 = (22'h93b !== 20'h10d4);
		#10; r150 = ( ( ^ ( r156)) && (((( ( | ( r211)) != r229) + (r249 - ((r17 ?  ( + (  ( ~ ( (( ( ! (  ( & ( 31'h6a65)))) || r174) && r229))))) : (r109 - r100)) | (((31'h15d == (12'h2b & ( ( ! ( r246)) + $time))) <= r14) >= ((30'h34b2 != r120) - (((((r100 === (r251 ^ 22'h665)) ? ((19'h2712 || r233) - ((8'h17 * 32'h4a8) * (12'h98c % 11'h480))) : r56) > (r104 ^ r14)) -  ( ~ (  ( - ( ( ( | ( (4'h2 !== 29'h34bc))) !=  ( & ( r57)))))))) >=  ( ^ ( r63)))))))) && 7'h66) !== 14'h1b9f));
		#10; r162 = r235;
		#10; r172 = (r216 > ($time > (28'h5158 % r196)));
		#10; r184 = (( ( - ( r45)) != (((r130 >=  ( ! ( (r19 === $stime)))) > (14'h520 /  ( ^ ( 15'h5fdb)))) && $time)) ===  ( & ( (r242 &&  ( ^ ( (((r120 * r148) <= ((r231 < r248) | r48)) != r187)))))));
		#10; r17 = 11'h50b;
		#10; r55 = (12'h425 !== $time);
		#10; r153 = r221;
		#10; r74 = 29'h4919;
		#10; r117 = r42;
		#10; r28 = $time;
		#10; r32 = (r204 ? ((r140 >= $time) > (r15 %  ( | ( ((9'h109 * r58) * r240))))) : ( ( & ( ((5'h8 / r5) ? 3'h2 : r72))) > (3'h0 -  ( ^ ( r104)))));
		#10; r11 = (r105 | ((r67 >= (((((11'h6cc == 20'h5279) - (((( ( ^ ( 2'h0)) >= (25'h262e % (((1'h1 ^ 4'h5) < (32'h34e3 + 32'h3f3f)) ^ r81))) !== (3'h1 - r162)) & ( ( + (  ( ! ( r171)))) === ((r95 && 3'h1) % 11'h241))) < $time)) / 14'h3e43) - r219) - 5'h0)) % ((22'h6f46 < ( ( ^ (  ( ! ( ((15'h4328 == (9'h7a < r234)) > r75))))) && r179)) &&  ( & ( (r174 * r120))))));
		#10; r152 = ( ( & ( r53)) % (r193 - ((((r106 % r173) && r85) / $time) *  ( - ( r82)))));
		#10; r181 = r166;
		#10; r189 = 23'h5062;
		#10; r129 = 12'h998;
		#10; r39 = 32'h51e9;
		#10; r16 = (($time % 12'h63f) + r134);
		#10; r223 = 12'h62;
		#10; r51 = (( ( ^ ( 9'h6b)) &  ( ! ( (28'h7eb0 | (r13 > (((r131 % (r176 != ((21'h7647 === ((22'h4cf1 ^ r217) * ( ( + ( 15'h40e1)) / r15))) ^ r191))) / ($stime || ( ( & ( ( ( - ( 7'h51)) <= ((19'h3479 > ((11'h518 > 25'h3c63) | (11'h243 ? 14'h3d56 : 11'h19e))) == (((25'h42 == 29'h4a37) > r19) * r255))))) && r196))) % r91)))))) + r104);
		#10; r177 = (22'h187d + (23'h2808 < ((r46 >=  ( - ( 8'hef))) & ((20'h68db !=  ( - ( r158))) + r185))));
		#10; r194 = $stime;
		#10; r219 = r208;
		#10; r94 = r73;
		#10; r61 = ((r25 - 26'h3cec) &&  ( - ( (r171 & r51))));
		#10; r249 = (17'h1cad > $stime);
		#10; r238 = (((r100 === r94) ? ((( ( + ( 31'h39d9)) == r226) === (r220 + $time)) ===  ( ^ ( ( ( ^ ( 20'h5654)) != ((r147 +  ( | ( r163))) - $stime))))) : ((28'ha75 >= (19'h59e0 - 32'h11eb)) > 25'h2ad6)) > 6'h32);
		#10; r176 = r71;
		#10; r239 =  ( & ( (r64 ?  ( - ( 25'h3d72)) : r249)));
		#10; r34 = ((((((r153 == r230) && (( ( ^ ( ((r127 != (((28'h4dc6 !=  ( ! (  ( ! ( 18'h3da9))))) -  ( ! ( ((9'h12e % 4'h0) <= (19'h2020 | 20'h2df2))))) & r166)) != 24'h3de8))) === (((r106 == ( ( & (  ( ~ ( r47)))) %  ( ~ ( ((r127 || r121) - (r238 !== (1'h1 >= 17'h5887))))))) -  ( & ( (12'h8b2 <= 17'hb10)))) +  ( + ( $time)))) ? 19'h55b5 :  ( | (  ( ^ (  ( ! ( (r147 ? (24'h3adc && 20'h2e20) : (r121 % ((( ( ~ ( 15'h1caa)) <= r178) <= (r238 ?  ( ! ( 27'h4907)) : (27'h1b95 && 19'h699e))) <= r225))))))))))) / r224) / r141) !=  ( + ( r154))) * (( ( ^ ( r176)) + 1'h0) || r214));
		#10; r195 = ( ( ! ( (20'h568d / ( ( | ( ( ( | ( (((r179 &&  ( ~ ( ( ( & ( ((14'h31b8 + 13'hab0) != 14'h758))) &  ( ! ( 4'h6)))))) < (11'h7d9 %  ( ! ( (21'h59ed != r91))))) - $stime))) + r10))) - r23)))) * 12'h86);
		#10; r198 = ((r185 == (24'h38c1 & (29'h636c !=  ( - ( (((r236 >=  ( & ( r244))) >= ( ( - ( ($time &  ( + ( r76))))) ? 17'h7d27 :  ( - ( 28'h42b0)))) -  ( + ( (19'hb62 === ((8'hc9 &&  ( ^ ( r143))) || (23'h13e0 !== (((17'h5c98 < r59) === (r141 >= ( ( ^ ( 27'h5389)) || (8'h5c != 10'h2ba)))) <= r136)))))))))))) < ((((23'h68e8 >= r212) ? (r115 < ( ( ^ (  ( ^ ( $stime)))) & (((((4'h7 ? ((r7 - $time) & (17'h6c4b > (26'h1d90 !== (22'h6c66 < 6'h2f)))) : 26'h1f77) >= (20'h5a16 >  ( ^ (  ( ^ ( ((11'h2f1 > 10'h3f7) ^  ( - ( 32'h719e))))))))) - $time) == 24'h11e0) * ( ( + ( r122)) - 5'h6)))) : r221) >=  ( | (  ( + ( (14'h2a24 - (16'h6dd0 >= 25'h1376))))))) > r54));
		#10; r79 = (( ( + ( ( ( + ( (((((20'h5369 && r249) ? (((r87 == (((5'h0 ? 14'h2f85 : 14'h1dae) / 30'h3c96) !== ((18'h7d54 >= 27'h19b) / (32'h6e73 != 32'h6d1e)))) === 15'h25af) *  ( + (  ( | ( (((24'h4069 !== 23'h5c26) && r36) &&  ( ! ( 29'h4aa6)))))))) : 9'h14e) / (9'h19b !== ( ( & ( $stime)) + 8'hb2))) || ((( ( | ( ((((26'h6ff8 ? 4'h9 : 10'h23d) ? (15'h1a1e || 17'h6cd9) : (11'h689 === 9'h1ac)) != 24'h16e8) == ( ( + ( r140)) & $time)))) & (30'h3029 > (4'ha * (r208 * ((8'h8b <= 27'h63d4) < r215))))) * (r123 > 3'h3)) | (27'h527f + r177))) + (19'h722e <= 6'h27)))) | (r183 >= ((7'h6a % ((10'h9e !== (r8 || ( ( ~ ( (r75 == (r104 !==  ( & ( 7'h23)))))) != ((r222 /  ( | ( 26'h1023))) !== $stime)))) > (r255 | $stime))) %  ( ! ( 23'h34ec))))))) == (( ( - ( 21'h6210)) * r195) !== ((28'h4979 > r232) | r22))) ^ (r125 * (r212 ^ (r10 != (((r201 >= 9'h39) < (( ( ~ ( (31'h2ca8 && ((18'h7958 - (((31'h50bf == 7'h73) === (10'h184 < 7'h0)) ||  ( & ( r100)))) + 17'h3580)))) >= ((r69 !== (r86 - (( ( & ( $time)) |  ( & (  ( - ( 22'h5f1b))))) >  ( ~ ( $time))))) ? 29'h6b06 : ((r236 >= 1'h1) < r25))) && 19'h2808)) === $time)))));
		#10; r100 = (((r202 <=  ( ~ ( r244))) == (r147 ? ( ( & ( (( ( | ( r167)) == r42) == r141))) + ( ( + (  ( + ( (((r254 ? $time : 18'h1c54) | r79) >= ((r25 === r206) != (r38 % r148))))))) * (7'h67 >= r127))) :  ( + ( ((( ( + ( (12'h4f9 !==  ( | ( r221))))) == ((r156 && (11'h216 | (((22'h66d5 || ((22'h1dd4 - 25'hd54) & (26'h133f | 12'h270))) * ( ( ! ( (23'h6438 > 6'h5))) ? ( ( - ( 7'h7b)) & r203) : ((23'h5cb4 ^ 28'h1157) <= (32'h4b39 + 23'h3ce5)))) <= (((30'h76b5 ? r69 : (24'h216b != 28'h41db)) |  ( + ( r123))) * ($stime !== ((28'hf8e >= 22'h7349) > r202)))))) ^ ((r9 != r99) ||  ( & ( (r224 >= r134)))))) || r56) ^ r235))))) ? r79 : ( ( ^ ( ((15'h2d1e !== ((((5'h11 >= $stime) | 6'h2a) * ((27'hfa0 <  ( ~ (  ( | (  ( ~ ( r156))))))) & (11'hb2 * r48))) === r166)) ==  ( + ( (((r136 ||  ( + ( ((( ( - ( 5'h1b)) == ( ( + ( (19'h2300 / 10'h2df))) <= 2'h0)) ^ ( ( ! (  ( - ( 10'hd2)))) / (((27'h3b64 * 16'h3f17) - (10'h3d4 | 5'h18)) == r74))) * r112)))) < 28'h4d35) *  ( | ( ( ( ! ( (29'h355f <=  ( ! ( r124))))) | ((r221 |  ( - ( ((r23 + r167) >  ( ! ( r106)))))) % r22)))))))))) ^  ( ! ( ((r246 & 27'h151c) >= 5'h1e)))));
		#10; r54 = 10'h1cf;
		#10; r51 = ((r132 >=  ( | ( (r228 && 24'h35b3)))) / 3'h7);
		#10; r43 = (r28 >  ( - ( (r24 % ((r100 & (r249 % r181)) ? 28'h6c6d : (26'h6a62 && (r47 > ((13'haae != (r63 ==  ( ! ( ((((r48 || 4'h4) ^ (r249 >= (18'h3348 ? 30'h2e36 : 23'hf79))) /  ( & ( r72))) ^ ((r147 || (r217 >= (29'h77b4 >= 14'h585))) >=  ( ^ ( 10'h1ba)))))))) % ((( ( + (  ( - ( $stime)))) | $stime) > 30'h2161) % ($time % (( ( ~ (  ( & ( 5'h3)))) == r206) || r203)))))))))));
		#10; r49 =  ( + ( (( ( ^ ( (32'h73e8 <= ((13'h372 < ((r196 /  ( ! ( ( ( - ( (r29 / (17'h609c && 6'h2f)))) / r103)))) && ((r245 + 21'h5feb) === (r195 < (r240 % ((((23'h27da + 26'hc96) ==  ( & ( 25'h7a84))) >= ( ( - ( 29'h33a4)) !== (5'he * 3'h0))) % (( ( + ( 1'h0)) ^ (18'h6e7e != 30'h3fba)) & $stime))))))) * 16'h88f)))) * 10'h3fb) < ((($stime % 26'h3cd3) * ((((r63 !== 32'h1ea4) + (13'hd6c != 3'h4)) < (($time > 31'h6440) + ((r51 && ( ( ! ( r108)) == (r28 % 10'h25e))) ^ r75))) - 22'h20d8)) & 10'h396))));
		#10; r248 = 23'h1af5;
		#10; r125 = 17'h1787;
		#10; r156 = $time;
		#10; r200 = (($stime ? 20'h295e : r19) != r135);
		#10; r209 = (( ( ~ ( (((((r97 + r9) - 12'h97a) - r11) > ((((r69 ==  ( ~ ( (r37 /  ( & ( (((26'h2658 == 3'h1) && (12'h375 && 11'h76f)) * r35))))))) != 10'h290) % (r169 &&  ( ! (  ( + ( (($time % (r31 % (r216 | (13'h4f9 * 11'hd9)))) / r216))))))) * r94)) / (r8 + r209)))) < 1'h0) >  ( | ( r166)));
		#10; r165 = (9'hd2 - r156);
		#10; r126 = 7'h15;
		#10; r90 = ((r171 != ( ( ~ ( ((((20'h4f9f <= (r116 & r103)) >= ((r111 % 15'h61e6) == r145)) == $stime) == 29'h475b))) &&  ( - ( (r207 ? r100 : ( ( - (  ( ! ( 9'hd0)))) /  ( | ( $time)))))))) / r85);
		#10; r82 = 26'h4010;
		#10; r112 = r191;
		#10; r222 = 9'h31;
		#10; r185 = (( ( ~ (  ( & ( ($stime != (( ( | ( (1'h1 ^ $time))) != r163) < (((r136 === (r43 % $stime)) == r192) <=  ( + ( (r211 ^ (20'h60aa !=  ( ^ ( (( ( ^ ( (4'h1 <= 20'h42af))) ?  ( ! ( (1'h1 - 16'h105))) : (16'h18a6 && 10'h379)) | r63)))))))))))))) && (r71 ^ 30'h3a7e)) >= r52);
		#10; r63 = (( ( ! ( 19'h71d2)) || r72) && r82);
		#10; r67 = r122;
		#10; r201 = (r110 ^  ( | ( ($stime ? ((r117 - 4'h5) && ( ( - ( (r35 / (18'h7494 == (22'h463d %  ( & ( 22'h302e))))))) / (r141 % ((4'h2 | (r78 * 19'h741d)) <=  ( + ( ($stime != 16'h441e))))))) : r252))));
		#10; r14 = 8'h25;
		#10; r227 = ( ( ! ( (((( ( ! ( (((12'ha44 - 13'h5b3) ? ((r235 || ((((8'he9 ? 27'h1dce : 10'h4a) !==  ( - ( 32'h4efe))) !== 24'h5642) > r86)) <= (7'h76 % ((((5'h1e | 28'h60ab) != (13'hd0a + 21'h76b8)) === ((19'h402 % 20'h77e0) || r205)) + r145))) : r242) ==  ( ! ( ( ( | (  ( | ( (r120 <= ( ( & ( 8'h25)) - $time)))))) >  ( | ( ( ( - ( r5)) ? 11'h276 : ( ( ^ ( 31'hbc7)) <= r90)))))))))) -  ( - ( (((( ( + ( r232)) && $stime) & $time) * r150) ? r41 :  ( | ( ((18'h22f3 / 4'h6) == (r76 ? ( ( | ( ($stime && (5'h18 <= 12'h483)))) & $stime) : ((((9'h54 <= 32'h2f44) | (3'h5 <= 16'h57af)) > 30'h3427) < $time))))))))) - (( ( | ( ( ( ~ (  ( ! ( ((r235 > r232) ^  ( ^ (  ( | (  ( - ( 3'h0))))))))))) && r240))) + r116) - ( ( ^ (  ( ! ( r19)))) % (r176 != r71)))) ? (r82 != 19'h5d16) : ((((r247 + (r124 - ((10'h13b > r155) === (r73 / $stime)))) < r246) / ((r9 - r190) + ((r25 ^ ((25'h720b / ( ( | ( ((19'h3f50 && 4'h8) & (30'h1773 || 5'h13)))) > (r150 | 19'h5393))) || ((r12 >= (((17'h434d === 8'hd9) * 29'h5a0b) > r21)) & r129))) * ( ( - ( r99)) == r227)))) < (22'h791f <= 5'h1b))) + r18))) && ((8'h71 == 3'h7) !== r85));
		#10; r112 = $stime;
		#10; r9 =  ( ^ ( (r91 !==  ( + ( ((r23 >= r175) | (((14'h144a + ((3'h6 * (r67 || ((( ( | ( (2'h2 != 22'h5093))) && 17'h18af) + (32'h3d27 > 9'h11)) - (((12'h474 && $time) != ((13'h1f06 * 4'he) == (6'h20 + 20'h106))) ?  ( ! (  ( & (  ( - ( 18'h7b24)))))) : r173)))) != 6'h15)) + 4'h1) & $time)))))));
		#10; r143 = 14'h2865;
		#10; r123 = 6'h3d;
		#10; r68 = (10'h296 *  ( ^ ( ( ( + ( ((((((26'h6a45 -  ( - ( ((27'h5a8b ^ (r216 || (19'h67a3 + 16'h4b36))) ^  ( + ( 2'h3)))))) && 14'h1816) || r144) *  ( - ( r153))) / r192) ^ ((r128 * r13) &  ( | ( r212)))))) != ((11'h5f0 ^ 9'h17e) == ((27'h62f3 > r48) | r84))))));
		#10; r233 = r38;
		#10; r11 = r39;
		#10; r138 = (( ( - ( 25'h745)) === (23'h560d >=  ( | (  ( ~ ( r208)))))) ^ (((r193 % r112) % (25'h2df3 === 30'h2e15)) || r198));
		#10; r122 = 24'h62ec;
		#10; r255 = 24'h4ba0;
		#10; r107 = (((r202 || ((19'h6de4 | 18'h4463) | (7'h7 + (2'h0 %  ( - (  ( ! ( ( ( ^ ( (r46 !== ((29'h1a74 ^ ( ( - ( 7'h69)) !=  ( ! ( 15'h777)))) - (((9'h90 / 29'h787c) && (29'h2626 !== 10'h11c)) | (5'hb ==  ( ! ( 14'h2aec)))))))) || r224))))))))) <= ((($stime % r96) || (( ( & ( ( ( ^ ( ((((((8'hc5 < 30'h3fbc) ? r59 : (26'h6bb6 !== 20'h4c53)) & ( ( ~ ( 32'h1e0d)) !=  ( - ( 14'h85c)))) !== ((r245 ? 18'h5cb8 : (6'h8 | 31'h321c)) != ((15'h260b - 18'h4db3) >= (18'h4dd >= 16'h703b)))) % r225) < r158))) + 22'h6c04))) >= (r216 + $time)) ? (((r243 |  ( ~ (  ( ^ ( 3'h4))))) < ((((26'h5eda ? $time : (r243 + 32'h15fb)) != 31'h1d73) < ((r52 <= r10) < (((31'h5a7c === (r163 & (10'h2e4 >= 29'h1549))) || r119) != ($time !== r184)))) ||  ( ^ ( ( ( ~ ( (((12'h669 ^ (25'h5139 | 22'h54d2)) & r123) !== 7'h56))) != r7))))) / (r81 | 8'h39)) :  ( ! ( r60)))) ?  ( ^ ( r135)) : r94)) / 21'h5e3f);
		#10; r80 = ((r16 ? r183 : ($time <= r178)) /  ( + ( ( ( | ( ((r54 !== r222) + (( ( ~ (  ( + ( 3'h3)))) && ((((((( ( ! ( 2'h1)) != (23'h4dc1 || 25'h6418)) & ((15'h3134 + 2'h1) * (4'h4 ? 29'h7aeb : 24'h1db3))) || r131) < r248) + ($time &  ( | ( r78)))) | ((((8'he9 || ((28'h64f2 != 31'h5ecb) == (5'h10 !== 16'h7020))) || (((20'h1b88 % 27'h7c75) - (1'h0 === 5'h0)) %  ( | ( (12'h4b9 & 19'h5c3b))))) - (17'he76 <= 2'h3)) /  ( ~ ( r73)))) <= (17'h386e | (r194 %  ( - (  ( ! ( ($time - r125))))))))) > 15'h7f04)))) === 13'h1828))));
		#10; r37 = (($stime == ((r41 !==  ( | ( 27'h1da6))) === (r35 ===  ( & ( 27'h2564))))) || ((16'h512e ? r184 : $stime) & 25'h56a4));
		#10; r96 =  ( - (  ( ~ ( r31))));
		#10; r246 = $stime;
		#10; r251 = 28'h62ae;
		#10; r143 = r4;
		#10; r123 = (r86 - $time);
		#10; r65 = r247;
		#10; r188 = r248;
		#10; r89 = ( ( & ( r73)) & r43);
		#10; r185 = 1'h1;
		#10; r45 = (( ( | (  ( ^ ( 24'h1a2d)))) !== r2) <=  ( + ( 22'h7447)));
		#10; r92 = (($stime %  ( ^ ( (((r236 ? (((((10'h240 ? 22'h7a0d : r163) * 20'h71a2) >= ( ( - ( r186)) < ((r104 * (((27'h7436 === 20'hbfb) || (13'h1d62 | 26'h6221)) != ((29'h823 && 6'h34) ^ r170))) % ( ( - ( r11)) % (((32'h611e / 31'h3c4c) +  ( & ( 20'h30a4))) - ((12'h85b == 26'hfd9) < 22'h74bb)))))) | (24'h4b4e >  ( ! (  ( | ( (( ( + ( (29'h63b9 >= 31'h5396))) < (28'h24a0 & (4'h5 | 6'h1c))) |  ( - ( ((13'h6a7 & 5'h3) >=  ( | ( 1'h0)))))))))))) % (r164 === r50)) : 13'h25d) == 19'h4390) || r105)))) | r180);
		#10; r23 = (5'h5 ^  ( ! ( $stime)));
		#10; r8 = ($time ? (32'h605f >= ((r233 >  ( ~ ( ( ( ^ ( (r28 * 26'h48ea))) ^ (((16'h617e & (10'he4 / r234)) ? 29'h1e10 : ( ( & ( 11'h22)) | $stime)) *  ( | (  ( - ( ((r200 | r159) == ((r226 < ((22'h50da ^ r22) >= (19'h5845 >  ( + ( 16'h3e29))))) !== (( ( ! ( (29'h34fe && 6'hc))) !== ((26'h35c4 < 20'h5230) * (30'h14f8 === 6'he))) < (((10'hc9 >= 12'h616) / (24'h6357 ^ 29'he15)) >= 31'h2b58))))))))))))) - ( ( ^ ( 10'h2af)) == ((32'h50d6 < 24'h30c0) > 22'h570e)))) : r232);
		#10; r245 = (r165 === (r147 === r18));
		#10; r57 =  ( - ( r200));
		#10; r208 =  ( | ( (r75 > 5'h2)));
		#10; r153 =  ( + ( r49));
		#10; r80 = ( ( - ( (r204 === ((4'h8 <= 14'h3eda) / r161)))) % ( ( | ( 17'h27bf)) != r40));
		#10; r230 = ((r196 & ((28'h44ec / r235) - ( ( | ( r84)) ^  ( | ( r199))))) & ( ( - ( (r215 % ((21'h63b8 < (r247 || ((9'h1b4 - 5'he) ? r129 : (((7'h48 / r63) < 30'h6df7) <= $time)))) - (r161 <= r141))))) == $time));
		#10; r58 = r227;
		$displayb("r0 = ",r0);
		$displayb("r1 = ",r1);
		$displayb("r2 = ",r2);
		$displayb("r3 = ",r3);
		$displayb("r4 = ",r4);
		$displayb("r5 = ",r5);
		$displayb("r6 = ",r6);
		$displayb("r7 = ",r7);
		$displayb("r8 = ",r8);
		$displayb("r9 = ",r9);
		$displayb("r10 = ",r10);
		$displayb("r11 = ",r11);
		$displayb("r12 = ",r12);
		$displayb("r13 = ",r13);
		$displayb("r14 = ",r14);
		$displayb("r15 = ",r15);
		$displayb("r16 = ",r16);
		$displayb("r17 = ",r17);
		$displayb("r18 = ",r18);
		$displayb("r19 = ",r19);
		$displayb("r20 = ",r20);
		$displayb("r21 = ",r21);
		$displayb("r22 = ",r22);
		$displayb("r23 = ",r23);
		$displayb("r24 = ",r24);
		$displayb("r25 = ",r25);
		$displayb("r26 = ",r26);
		$displayb("r27 = ",r27);
		$displayb("r28 = ",r28);
		$displayb("r29 = ",r29);
		$displayb("r30 = ",r30);
		$displayb("r31 = ",r31);
		$displayb("r32 = ",r32);
		$displayb("r33 = ",r33);
		$displayb("r34 = ",r34);
		$displayb("r35 = ",r35);
		$displayb("r36 = ",r36);
		$displayb("r37 = ",r37);
		$displayb("r38 = ",r38);
		$displayb("r39 = ",r39);
		$displayb("r40 = ",r40);
		$displayb("r41 = ",r41);
		$displayb("r42 = ",r42);
		$displayb("r43 = ",r43);
		$displayb("r44 = ",r44);
		$displayb("r45 = ",r45);
		$displayb("r46 = ",r46);
		$displayb("r47 = ",r47);
		$displayb("r48 = ",r48);
		$displayb("r49 = ",r49);
		$displayb("r50 = ",r50);
		$displayb("r51 = ",r51);
		$displayb("r52 = ",r52);
		$displayb("r53 = ",r53);
		$displayb("r54 = ",r54);
		$displayb("r55 = ",r55);
		$displayb("r56 = ",r56);
		$displayb("r57 = ",r57);
		$displayb("r58 = ",r58);
		$displayb("r59 = ",r59);
		$displayb("r60 = ",r60);
		$displayb("r61 = ",r61);
		$displayb("r62 = ",r62);
		$displayb("r63 = ",r63);
		$displayb("r64 = ",r64);
		$displayb("r65 = ",r65);
		$displayb("r66 = ",r66);
		$displayb("r67 = ",r67);
		$displayb("r68 = ",r68);
		$displayb("r69 = ",r69);
		$displayb("r70 = ",r70);
		$displayb("r71 = ",r71);
		$displayb("r72 = ",r72);
		$displayb("r73 = ",r73);
		$displayb("r74 = ",r74);
		$displayb("r75 = ",r75);
		$displayb("r76 = ",r76);
		$displayb("r77 = ",r77);
		$displayb("r78 = ",r78);
		$displayb("r79 = ",r79);
		$displayb("r80 = ",r80);
		$displayb("r81 = ",r81);
		$displayb("r82 = ",r82);
		$displayb("r83 = ",r83);
		$displayb("r84 = ",r84);
		$displayb("r85 = ",r85);
		$displayb("r86 = ",r86);
		$displayb("r87 = ",r87);
		$displayb("r88 = ",r88);
		$displayb("r89 = ",r89);
		$displayb("r90 = ",r90);
		$displayb("r91 = ",r91);
		$displayb("r92 = ",r92);
		$displayb("r93 = ",r93);
		$displayb("r94 = ",r94);
		$displayb("r95 = ",r95);
		$displayb("r96 = ",r96);
		$displayb("r97 = ",r97);
		$displayb("r98 = ",r98);
		$displayb("r99 = ",r99);
		$displayb("r100 = ",r100);
		$displayb("r101 = ",r101);
		$displayb("r102 = ",r102);
		$displayb("r103 = ",r103);
		$displayb("r104 = ",r104);
		$displayb("r105 = ",r105);
		$displayb("r106 = ",r106);
		$displayb("r107 = ",r107);
		$displayb("r108 = ",r108);
		$displayb("r109 = ",r109);
		$displayb("r110 = ",r110);
		$displayb("r111 = ",r111);
		$displayb("r112 = ",r112);
		$displayb("r113 = ",r113);
		$displayb("r114 = ",r114);
		$displayb("r115 = ",r115);
		$displayb("r116 = ",r116);
		$displayb("r117 = ",r117);
		$displayb("r118 = ",r118);
		$displayb("r119 = ",r119);
		$displayb("r120 = ",r120);
		$displayb("r121 = ",r121);
		$displayb("r122 = ",r122);
		$displayb("r123 = ",r123);
		$displayb("r124 = ",r124);
		$displayb("r125 = ",r125);
		$displayb("r126 = ",r126);
		$displayb("r127 = ",r127);
		$displayb("r128 = ",r128);
		$displayb("r129 = ",r129);
		$displayb("r130 = ",r130);
		$displayb("r131 = ",r131);
		$displayb("r132 = ",r132);
		$displayb("r133 = ",r133);
		$displayb("r134 = ",r134);
		$displayb("r135 = ",r135);
		$displayb("r136 = ",r136);
		$displayb("r137 = ",r137);
		$displayb("r138 = ",r138);
		$displayb("r139 = ",r139);
		$displayb("r140 = ",r140);
		$displayb("r141 = ",r141);
		$displayb("r142 = ",r142);
		$displayb("r143 = ",r143);
		$displayb("r144 = ",r144);
		$displayb("r145 = ",r145);
		$displayb("r146 = ",r146);
		$displayb("r147 = ",r147);
		$displayb("r148 = ",r148);
		$displayb("r149 = ",r149);
		$displayb("r150 = ",r150);
		$displayb("r151 = ",r151);
		$displayb("r152 = ",r152);
		$displayb("r153 = ",r153);
		$displayb("r154 = ",r154);
		$displayb("r155 = ",r155);
		$displayb("r156 = ",r156);
		$displayb("r157 = ",r157);
		$displayb("r158 = ",r158);
		$displayb("r159 = ",r159);
		$displayb("r160 = ",r160);
		$displayb("r161 = ",r161);
		$displayb("r162 = ",r162);
		$displayb("r163 = ",r163);
		$displayb("r164 = ",r164);
		$displayb("r165 = ",r165);
		$displayb("r166 = ",r166);
		$displayb("r167 = ",r167);
		$displayb("r168 = ",r168);
		$displayb("r169 = ",r169);
		$displayb("r170 = ",r170);
		$displayb("r171 = ",r171);
		$displayb("r172 = ",r172);
		$displayb("r173 = ",r173);
		$displayb("r174 = ",r174);
		$displayb("r175 = ",r175);
		$displayb("r176 = ",r176);
		$displayb("r177 = ",r177);
		$displayb("r178 = ",r178);
		$displayb("r179 = ",r179);
		$displayb("r180 = ",r180);
		$displayb("r181 = ",r181);
		$displayb("r182 = ",r182);
		$displayb("r183 = ",r183);
		$displayb("r184 = ",r184);
		$displayb("r185 = ",r185);
		$displayb("r186 = ",r186);
		$displayb("r187 = ",r187);
		$displayb("r188 = ",r188);
		$displayb("r189 = ",r189);
		$displayb("r190 = ",r190);
		$displayb("r191 = ",r191);
		$displayb("r192 = ",r192);
		$displayb("r193 = ",r193);
		$displayb("r194 = ",r194);
		$displayb("r195 = ",r195);
		$displayb("r196 = ",r196);
		$displayb("r197 = ",r197);
		$displayb("r198 = ",r198);
		$displayb("r199 = ",r199);
		$displayb("r200 = ",r200);
		$displayb("r201 = ",r201);
		$displayb("r202 = ",r202);
		$displayb("r203 = ",r203);
		$displayb("r204 = ",r204);
		$displayb("r205 = ",r205);
		$displayb("r206 = ",r206);
		$displayb("r207 = ",r207);
		$displayb("r208 = ",r208);
		$displayb("r209 = ",r209);
		$displayb("r210 = ",r210);
		$displayb("r211 = ",r211);
		$displayb("r212 = ",r212);
		$displayb("r213 = ",r213);
		$displayb("r214 = ",r214);
		$displayb("r215 = ",r215);
		$displayb("r216 = ",r216);
		$displayb("r217 = ",r217);
		$displayb("r218 = ",r218);
		$displayb("r219 = ",r219);
		$displayb("r220 = ",r220);
		$displayb("r221 = ",r221);
		$displayb("r222 = ",r222);
		$displayb("r223 = ",r223);
		$displayb("r224 = ",r224);
		$displayb("r225 = ",r225);
		$displayb("r226 = ",r226);
		$displayb("r227 = ",r227);
		$displayb("r228 = ",r228);
		$displayb("r229 = ",r229);
		$displayb("r230 = ",r230);
		$displayb("r231 = ",r231);
		$displayb("r232 = ",r232);
		$displayb("r233 = ",r233);
		$displayb("r234 = ",r234);
		$displayb("r235 = ",r235);
		$displayb("r236 = ",r236);
		$displayb("r237 = ",r237);
		$displayb("r238 = ",r238);
		$displayb("r239 = ",r239);
		$displayb("r240 = ",r240);
		$displayb("r241 = ",r241);
		$displayb("r242 = ",r242);
		$displayb("r243 = ",r243);
		$displayb("r244 = ",r244);
		$displayb("r245 = ",r245);
		$displayb("r246 = ",r246);
		$displayb("r247 = ",r247);
		$displayb("r248 = ",r248);
		$displayb("r249 = ",r249);
		$displayb("r250 = ",r250);
		$displayb("r251 = ",r251);
		$displayb("r252 = ",r252);
		$displayb("r253 = ",r253);
		$displayb("r254 = ",r254);
		$finish(0);
	end
endmodule
