//
// Copyright (c) 2000 Paul Campbell (paul@verifarm.com)
//
//    This source code is free software; you can redistribute it
//    and/or modify it in source code form under the terms of the GNU
//    General Public License as published by the Free Software
//    Foundation; either version 2 of the License, or (at your option)
//    any later version.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program; if not, write to the Free Software
//    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
//
module compl1001;
	reg	[104:86]r0;
	reg	[261:230]r1;
	reg	[101:78]r2;
	reg	[216:215]r3;
	reg	[140:123]r4;
	reg	[70:53]r5;
	reg	[150:150]r6;
	reg	[143:133]r7;
	reg	[261:239]r8;
	reg	[228:211]r9;
	reg	[273:244]r10;
	reg	[42:21]r11;
	reg	[137:130]r12;
	reg	[103:96]r13;
	reg	[257:239]r14;
	reg	[230:205]r15;
	reg	[216:212]r16;
	reg	[64:40]r17;
	reg	[156:155]r18;
	reg	[103:94]r19;
	reg	[216:204]r20;
	reg	[170:165]r21;
	reg	[25:22]r22;
	reg	[125:105]r23;
	reg	[57:32]r24;
	reg	[261:250]r25;
	reg	[32:13]r26;
	reg	[251:246]r27;
	reg	[210:209]r28;
	reg	[121:119]r29;
	reg	[57:55]r30;
	reg	[255:253]r31;
	reg	[196:174]r32;
	reg	[26:26]r33;
	reg	[216:215]r34;
	reg	[238:224]r35;
	reg	[212:207]r36;
	reg	[32:11]r37;
	reg	[89:60]r38;
	reg	[246:237]r39;
	reg	[50:25]r40;
	reg	[43:29]r41;
	reg	[94:66]r42;
	reg	[235:222]r43;
	reg	[213:190]r44;
	reg	[102:81]r45;
	reg	[211:208]r46;
	reg	[108:91]r47;
	reg	[189:188]r48;
	reg	[97:84]r49;
	reg	[108:90]r50;
	reg	[124:116]r51;
	reg	[113:92]r52;
	reg	[278:254]r53;
	reg	[98:94]r54;
	reg	[43:42]r55;
	reg	[191:178]r56;
	reg	[230:211]r57;
	reg	[250:233]r58;
	reg	[236:229]r59;
	reg	[65:34]r60;
	reg	[155:132]r61;
	reg	[32:18]r62;
	reg	[253:253]r63;
	reg	[243:215]r64;
	reg	[133:109]r65;
	reg	[133:124]r66;
	reg	[66:51]r67;
	reg	[94:75]r68;
	reg	[31:23]r69;
	reg	[230:214]r70;
	reg	[75:55]r71;
	reg	[209:196]r72;
	reg	[200:181]r73;
	reg	[101:92]r74;
	reg	[43:34]r75;
	reg	[228:211]r76;
	reg	[171:169]r77;
	reg	[112:86]r78;
	reg	[257:252]r79;
	reg	[214:214]r80;
	reg	[279:254]r81;
	reg	[149:149]r82;
	reg	[80:53]r83;
	reg	[140:117]r84;
	reg	[265:238]r85;
	reg	[277:251]r86;
	reg	[71:45]r87;
	reg	[56:38]r88;
	reg	[95:91]r89;
	reg	[271:242]r90;
	reg	[187:174]r91;
	reg	[176:171]r92;
	reg	[100:88]r93;
	reg	[273:242]r94;
	reg	[137:111]r95;
	reg	[148:144]r96;
	reg	[168:159]r97;
	reg	[269:254]r98;
	reg	[149:145]r99;
	reg	[202:176]r100;
	reg	[37:26]r101;
	reg	[62:37]r102;
	reg	[47:36]r103;
	reg	[195:176]r104;
	reg	[124:93]r105;
	reg	[8:4]r106;
	reg	[170:161]r107;
	reg	[150:129]r108;
	reg	[54:40]r109;
	reg	[86:64]r110;
	reg	[132:111]r111;
	reg	[224:224]r112;
	reg	[262:232]r113;
	reg	[27:14]r114;
	reg	[99:97]r115;
	reg	[234:214]r116;
	reg	[66:52]r117;
	reg	[178:173]r118;
	reg	[83:52]r119;
	reg	[67:58]r120;
	reg	[110:82]r121;
	reg	[255:232]r122;
	reg	[41:19]r123;
	reg	[67:45]r124;
	reg	[179:178]r125;
	reg	[173:151]r126;
	reg	[35:20]r127;
	reg	[168:155]r128;
	reg	[129:112]r129;
	reg	[47:29]r130;
	reg	[199:186]r131;
	reg	[217:190]r132;
	reg	[241:212]r133;
	reg	[256:233]r134;
	reg	[129:116]r135;
	reg	[168:157]r136;
	reg	[230:211]r137;
	reg	[261:248]r138;
	reg	[39:27]r139;
	reg	[137:135]r140;
	reg	[169:142]r141;
	reg	[103:79]r142;
	reg	[118:118]r143;
	reg	[156:154]r144;
	reg	[234:208]r145;
	reg	[154:131]r146;
	reg	[211:183]r147;
	reg	[74:65]r148;
	reg	[161:145]r149;
	reg	[58:51]r150;
	reg	[268:253]r151;
	reg	[193:175]r152;
	reg	[148:120]r153;
	reg	[169:138]r154;
	reg	[213:210]r155;
	reg	[119:103]r156;
	reg	[104:83]r157;
	reg	[212:193]r158;
	reg	[172:172]r159;
	reg	[206:182]r160;
	reg	[176:159]r161;
	reg	[172:153]r162;
	reg	[119:110]r163;
	reg	[75:53]r164;
	reg	[5:5]r165;
	reg	[238:226]r166;
	reg	[258:230]r167;
	reg	[95:74]r168;
	reg	[231:216]r169;
	reg	[252:248]r170;
	reg	[98:79]r171;
	reg	[191:166]r172;
	reg	[161:154]r173;
	reg	[67:67]r174;
	reg	[214:207]r175;
	reg	[204:198]r176;
	reg	[131:118]r177;
	reg	[212:181]r178;
	reg	[258:248]r179;
	reg	[141:116]r180;
	reg	[201:198]r181;
	reg	[108:78]r182;
	reg	[83:72]r183;
	reg	[81:69]r184;
	reg	[144:140]r185;
	reg	[174:154]r186;
	reg	[191:171]r187;
	reg	[48:27]r188;
	reg	[260:251]r189;
	reg	[69:47]r190;
	reg	[259:246]r191;
	reg	[167:162]r192;
	reg	[245:237]r193;
	reg	[67:49]r194;
	reg	[133:108]r195;
	reg	[224:213]r196;
	reg	[126:108]r197;
	reg	[230:208]r198;
	reg	[80:59]r199;
	reg	[136:120]r200;
	reg	[62:44]r201;
	reg	[206:198]r202;
	reg	[284:254]r203;
	reg	[184:158]r204;
	reg	[32:13]r205;
	reg	[233:220]r206;
	reg	[69:59]r207;
	reg	[46:34]r208;
	reg	[181:156]r209;
	reg	[105:100]r210;
	reg	[240:228]r211;
	reg	[51:48]r212;
	reg	[149:144]r213;
	reg	[201:190]r214;
	reg	[234:215]r215;
	reg	[212:188]r216;
	reg	[98:79]r217;
	reg	[237:214]r218;
	reg	[105:96]r219;
	reg	[10:7]r220;
	reg	[134:105]r221;
	reg	[192:162]r222;
	reg	[202:180]r223;
	reg	[50:31]r224;
	reg	[50:26]r225;
	reg	[181:166]r226;
	reg	[146:117]r227;
	reg	[118:93]r228;
	reg	[222:202]r229;
	reg	[135:114]r230;
	reg	[78:51]r231;
	reg	[260:231]r232;
	reg	[172:142]r233;
	reg	[58:32]r234;
	reg	[245:232]r235;
	reg	[51:46]r236;
	reg	[198:167]r237;
	reg	[217:217]r238;
	reg	[130:121]r239;
	reg	[130:111]r240;
	reg	[28:0]r241;
	reg	[87:79]r242;
	reg	[60:58]r243;
	reg	[59:53]r244;
	reg	[200:178]r245;
	reg	[81:67]r246;
	reg	[110:104]r247;
	reg	[233:211]r248;
	reg	[139:129]r249;
	reg	[262:254]r250;
	reg	[177:175]r251;
	reg	[262:236]r252;
	reg	[111:94]r253;
	reg	[230:218]r254;
	reg	[191:164]r255;
	initial begin
		r0 = 32'h2eec;
		r1 = 32'h1584;
		r2 = 32'h47e5;
		r3 = 32'h587f;
		r4 = 32'hab8;
		r5 = 32'h71e9;
		r6 = 32'h4e49;
		r7 = 32'h6794;
		r8 = 32'h5c8e;
		r9 = 32'h1a61;
		r10 = 32'h55df;
		r11 = 32'h2da5;
		r12 = 32'h3d89;
		r13 = 32'h76ab;
		r14 = 32'h6d8e;
		r15 = 32'h66ed;
		r16 = 32'hc57;
		r17 = 32'h615c;
		r18 = 32'h29c0;
		r19 = 32'h7ed1;
		r20 = 32'h11c7;
		r21 = 32'h5f7a;
		r22 = 32'h59cc;
		r23 = 32'h36df;
		r24 = 32'h6217;
		r25 = 32'h35da;
		r26 = 32'h2827;
		r27 = 32'h418b;
		r28 = 32'h6fb;
		r29 = 32'h7839;
		r30 = 32'h114b;
		r31 = 32'h4ca3;
		r32 = 32'h3e6d;
		r33 = 32'h6e1d;
		r34 = 32'h5d63;
		r35 = 32'h3797;
		r36 = 32'h5a38;
		r37 = 32'h6969;
		r38 = 32'h8bb;
		r39 = 32'h716b;
		r40 = 32'hc42;
		r41 = 32'h6ac3;
		r42 = 32'h46ea;
		r43 = 32'h3a78;
		r44 = 32'h2b9c;
		r45 = 32'h2fa6;
		r46 = 32'hcbc;
		r47 = 32'h45e6;
		r48 = 32'h3e4b;
		r49 = 32'h646;
		r50 = 32'h4ce2;
		r51 = 32'h76e9;
		r52 = 32'h53d4;
		r53 = 32'h327;
		r54 = 32'h5359;
		r55 = 32'h35be;
		r56 = 32'h7c89;
		r57 = 32'h747c;
		r58 = 32'h6b9a;
		r59 = 32'h1864;
		r60 = 32'h6996;
		r61 = 32'h2f40;
		r62 = 32'h3d86;
		r63 = 32'h5b1b;
		r64 = 32'h1ca;
		r65 = 32'h1216;
		r66 = 32'hd10;
		r67 = 32'h649e;
		r68 = 32'h7727;
		r69 = 32'h59e1;
		r70 = 32'h48a8;
		r71 = 32'h521f;
		r72 = 32'h2928;
		r73 = 32'h2423;
		r74 = 32'h126b;
		r75 = 32'h4707;
		r76 = 32'h5fd4;
		r77 = 32'h3b16;
		r78 = 32'h300c;
		r79 = 32'h7c6a;
		r80 = 32'h2b87;
		r81 = 32'h78c;
		r82 = 32'hd80;
		r83 = 32'h4c4c;
		r84 = 32'h757b;
		r85 = 32'h4487;
		r86 = 32'h3e6c;
		r87 = 32'h3496;
		r88 = 32'hd19;
		r89 = 32'h5098;
		r90 = 32'h2a4f;
		r91 = 32'hdd6;
		r92 = 32'h3e02;
		r93 = 32'h38f8;
		r94 = 32'h4f6f;
		r95 = 32'h71ba;
		r96 = 32'h3adc;
		r97 = 32'h5a68;
		r98 = 32'h4884;
		r99 = 32'hd4a;
		r100 = 32'h68dd;
		r101 = 32'h33c8;
		r102 = 32'h127;
		r103 = 32'h5ae8;
		r104 = 32'h5818;
		r105 = 32'h4679;
		r106 = 32'h44f9;
		r107 = 32'h9;
		r108 = 32'h748a;
		r109 = 32'h2074;
		r110 = 32'h1593;
		r111 = 32'h4ab1;
		r112 = 32'h3be4;
		r113 = 32'h6c27;
		r114 = 32'h7331;
		r115 = 32'hab0;
		r116 = 32'h416;
		r117 = 32'h2213;
		r118 = 32'h41d;
		r119 = 32'h429e;
		r120 = 32'h1ea0;
		r121 = 32'h3827;
		r122 = 32'h46dd;
		r123 = 32'h6c97;
		r124 = 32'h6497;
		r125 = 32'h6ada;
		r126 = 32'h3b1c;
		r127 = 32'h4eb7;
		r128 = 32'h7779;
		r129 = 32'h7c0a;
		r130 = 32'h2d59;
		r131 = 32'h1b54;
		r132 = 32'h42b2;
		r133 = 32'h397;
		r134 = 32'h1151;
		r135 = 32'h58fe;
		r136 = 32'h9ea;
		r137 = 32'h2dbe;
		r138 = 32'h172d;
		r139 = 32'h4e38;
		r140 = 32'h1015;
		r141 = 32'h337;
		r142 = 32'h676c;
		r143 = 32'h6cf3;
		r144 = 32'h2338;
		r145 = 32'h170f;
		r146 = 32'h318e;
		r147 = 32'h79ce;
		r148 = 32'h18fc;
		r149 = 32'h3643;
		r150 = 32'h7986;
		r151 = 32'h6b10;
		r152 = 32'h7f4;
		r153 = 32'h7520;
		r154 = 32'h4fdd;
		r155 = 32'h3b61;
		r156 = 32'h49ae;
		r157 = 32'h365d;
		r158 = 32'h60a6;
		r159 = 32'h2c4b;
		r160 = 32'h117b;
		r161 = 32'h7f4;
		r162 = 32'h525;
		r163 = 32'h3475;
		r164 = 32'h23fe;
		r165 = 32'h71c5;
		r166 = 32'h443e;
		r167 = 32'h1599;
		r168 = 32'h7b77;
		r169 = 32'h11ea;
		r170 = 32'h6d9f;
		r171 = 32'h564a;
		r172 = 32'h64cd;
		r173 = 32'h22d8;
		r174 = 32'h3bad;
		r175 = 32'h1b68;
		r176 = 32'h615d;
		r177 = 32'h473a;
		r178 = 32'h282f;
		r179 = 32'h1d5e;
		r180 = 32'h5985;
		r181 = 32'h378d;
		r182 = 32'h5fbd;
		r183 = 32'h3522;
		r184 = 32'h6bef;
		r185 = 32'h2d7c;
		r186 = 32'h7fe6;
		r187 = 32'h3cea;
		r188 = 32'h659d;
		r189 = 32'h28f9;
		r190 = 32'hc24;
		r191 = 32'h40af;
		r192 = 32'h2eb9;
		r193 = 32'h6b1f;
		r194 = 32'h4581;
		r195 = 32'h3a63;
		r196 = 32'h381a;
		r197 = 32'h42cb;
		r198 = 32'h5105;
		r199 = 32'h55f1;
		r200 = 32'h3596;
		r201 = 32'h6f4;
		r202 = 32'h58e6;
		r203 = 32'h78f8;
		r204 = 32'h310a;
		r205 = 32'h5ace;
		r206 = 32'h146f;
		r207 = 32'ha48;
		r208 = 32'h422a;
		r209 = 32'h17a3;
		r210 = 32'h62ac;
		r211 = 32'h3518;
		r212 = 32'h7709;
		r213 = 32'h786c;
		r214 = 32'h63db;
		r215 = 32'h240d;
		r216 = 32'h3967;
		r217 = 32'h6332;
		r218 = 32'h3d92;
		r219 = 32'h6fec;
		r220 = 32'h3cbe;
		r221 = 32'h6c27;
		r222 = 32'h75af;
		r223 = 32'h3e19;
		r224 = 32'h410b;
		r225 = 32'h6e83;
		r226 = 32'h1004;
		r227 = 32'h4ad7;
		r228 = 32'h365d;
		r229 = 32'h5720;
		r230 = 32'h5abf;
		r231 = 32'h5b3e;
		r232 = 32'hd1f;
		r233 = 32'h7cd4;
		r234 = 32'h159b;
		r235 = 32'h52fb;
		r236 = 32'h3f25;
		r237 = 32'h2292;
		r238 = 32'h5fc9;
		r239 = 32'h69ca;
		r240 = 32'h5d77;
		r241 = 32'h7f3f;
		r242 = 32'h189c;
		r243 = 32'h3cb5;
		r244 = 32'h2ee1;
		r245 = 32'h6755;
		r246 = 32'h1ef7;
		r247 = 32'h370a;
		r248 = 32'h2b36;
		r249 = 32'h743a;
		r250 = 32'h1b77;
		r251 = 32'hf1d;
		r252 = 32'h5f68;
		r253 = 32'h455e;
		r254 = 32'h415f;
		r255 = 32'h52c2;
		#10; r73 = r189;
		#10; r132 = 11'h783;
		#10; r86 = ( ( & ( (14'h1136 ^ ((25'hd6c == $time) * r2)))) != 26'h1ef2);
		#10; r246 =  ( | ( 22'h6337));
		#10; r35 = (r155 * ((r190 > (((((((r127 %  ( | ( r81))) & r150) | r11) !== (((r207 <= (22'h4d2b ? ((r158 ==  ( - ( r219))) | 13'hdae) : r43)) != ((r97 > ((r240 != ((26'h259a * 13'h465) >= (5'h2 * 11'h7ed))) % (((12'h279 < 28'h3026) || 4'h1) && r111))) &  ( ! (  ( ! ( (16'h7a99 <= 4'h6))))))) & 26'h5fa4)) && (((r15 | (( ( | (  ( ~ ( (r235 && 31'h2eeb))))) / r90) !== r56)) <= ((22'h640f !== r182) <= (31'h1b37 !== ( ( | ( (((9'hc9 / 32'h7c3b) - (8'ha6 - 3'h2)) == ((12'h36b - 9'h171) <  ( + ( 23'h425)))))) % r72)))) + $time)) > r1) !== 18'h6d7b)) >= 28'h6e25));
		#10; r144 = 4'h9;
		#10; r206 = ( ( | ( 12'h4ff)) | 17'h43ef);
		#10; r138 = $time;
		#10; r74 = 22'h38ad;
		#10; r49 = r2;
		#10; r50 = ((31'h744c ? ((r164 && r191) >= 16'h6c50) : ((r137 / ((1'h0 ^ ((r169 >= (((20'h5ab3 ==  ( & (  ( & ( (21'hb12 < (7'h16 || 10'h24e))))))) != r155) -  ( | (  ( + ( ( ( ! ( r166)) % (26'h296c > 32'h62ed)))))))) ===  ( + (  ( | ( r187)))))) - r92)) * r99)) >= r189);
		#10; r150 = ((12'h24d != r248) /  ( & ( (((r34 -  ( ! ( 20'h40cd))) === (((7'h52 > (25'h7f1d || 1'h1)) && 5'h12) ?  ( ^ ( (r61 &&  ( ~ ( ( ( + (  ( ! ( (r73 <=  ( | ( ( ( & ( 28'h57c)) / (24'h60a8 < 28'h7acc))))))))) | (8'h61 <  ( ! ( (r184 ===  ( ~ ( (r72 == (15'h508 / 24'h5073)))))))))))))) : r24)) | r86))));
		#10; r73 = ( ( + ( ( ( ~ ( ((((20'h23e2 === ((11'h649 ^ 21'hfee) | ((r35 % 30'h856) <= r67))) !== ((r183 || (((r19 / (15'h304d + 25'h523a)) && 17'h7692) - r178)) - (((((25'h34f5 || r199) === r255) <= r12) !== (((((5'hb / 5'h11) == (5'h17 | 24'h408)) / (r255 ^ r181)) &&  ( & ( 14'h2e37))) === ((17'h1e79 <= r84) / (r0 !==  ( ^ ( (26'h587b <= 20'h7403))))))) >=  ( - ( r184))))) !==  ( - ( r248))) === $time))) * 12'h5))) || r191);
		#10; r134 = (1'h1 === 24'h12a0);
		#10; r214 = 30'h3839;
		#10; r255 = 30'h242b;
		#10; r7 = 9'h132;
		#10; r130 = r65;
		#10; r64 = r162;
		#10; r174 = ((r91 <= (r231 +  ( - ( 1'h1)))) <= ((((r93 <= (r183 / ( ( & (  ( ^ (  ( ^ ( 1'h1)))))) <= r75))) * 12'ha95) & r27) | ((((((20'hf1f === ((r175 >= 20'h3632) | ((r109 & (r88 < r248)) < 10'h2e5))) & r37) % $stime) || ( ( + (  ( ! ( r160)))) & r17)) > ( ( | ( (r124 &  ( - (  ( - ( (22'hd2b !=  ( ! ( r196)))))))))) && r84)) | (r51 / 16'h5f0d))));
		#10; r41 = ( ( ^ ( ( ( ^ ( ((3'h6 >= (r215 & (31'h3d8b &&  ( ^ ( 5'h11))))) <= $time))) &  ( & ( r7))))) * ( ( - ( (12'he7e ?  ( + ( ((3'h2 ^ r250) & (r214 <= (r19 - r249))))) : (r140 | r104)))) || r250));
		#10; r195 = 9'h1ac;
		#10; r242 = 21'h527c;
		#10; r143 = ((((((r68 ? (6'h1e ?  ( ^ ( 26'h4f04)) :  ( - ( ( ( - ( $time)) - (( ( + ( r96)) !== (r185 / 6'h22)) ? r133 : r2))))) : r20) * ((28'h20ec % r109) /  ( + ( ( ( & ( 1'h0)) | (13'h13f1 === ((r96 - r204) *  ( | ( 1'h0))))))))) === ((23'h4c6b / (20'h7a3b === r184)) == (( ( ! ( ( ( + ( (((7'h59 ? ((3'h4 <= 13'had1) | 15'h1a5c) : r123) % $stime) ==  ( + ( (((15'h74fe === 2'h0) ==  ( + ( 3'h0))) <= ((26'h2e1 | 8'h3b) + (16'h76a4 == 26'h645a)))))))) +  ( + ( ((r123 & (r37 != (r211 >= (21'hcee < 18'h2845)))) >= (27'h5efd ^ r116))))))) | ((25'h4cd6 + r74) ? r115 : ((r133 - ((r198 ? r55 : (($stime % 17'h38a5) | $time)) ===  ( ~ ( r217)))) ? (r250 !== 19'h49e1) :  ( ! ( r15))))) == r224))) - ((r244 > (r229 -  ( & ( (( ( + ( r244)) !=  ( ! ( ((29'h6d1b === 10'h364) - ((17'h43c9 &  ( + ( r238))) == r113))))) % 30'h7539))))) &  ( | ( 23'h4205)))) | 5'h19) <=  ( ! ( r92)));
		#10; r74 = r232;
		#10; r31 = ( ( ~ ( r181)) &&  ( - ( 7'h8)));
		#10; r75 = (6'h10 === r188);
		#10; r75 = ( ( & ( $stime)) +  ( - ( ((( ( | ( (16'h1c8a % 32'h503f))) ? ((r161 ^ r59) ==  ( ! (  ( - ( (((r191 === r182) == ( ( + (  ( | ( r168)))) > ( ( | ( 1'h1)) * (( ( ^ ( 32'h2923)) != (14'h3cd7 * 24'h1162)) > (25'h7bc2 - 6'hd))))) - r31)))))) : ((4'hd &  ( ^ ( (r130 - ((r96 === r154) == (32'h2fba >=  ( | ( 4'h3)))))))) >=  ( & ( (((r253 !== 18'h4189) >= (11'h679 < r133)) * r109))))) != $time) !== ( ( ~ ( (((21'h5dd3 / (10'h22e ^ (( ( ! (  ( + (  ( & ( (21'h5c32 * 12'h7e))))))) - ((((16'h132e || 23'hf58) <= 21'h1302) ^ ((2'h1 | 4'hb) - r113)) & (r207 || 24'h1190))) || ((r224 && r246) > 7'h19)))) % ( ( ~ ( r150)) - ((1'h1 & 24'h7aa2) | ($stime !== r24)))) >= 14'h29de))) !==  ( + ( 10'h207)))))));
		#10; r195 = 4'h7;
		#10; r129 = r208;
		#10; r152 = r144;
		#10; r9 = (( ( ! (  ( & ( (r39 >= r176))))) - 5'h6) ^ 12'h837);
		#10; r159 =  ( + ( ((r132 <= (((( ( + ( (24'h5c17 + r12))) == 24'h3ca7) > r164) >= ( ( ^ ( r114)) > r126)) < ((r0 &  ( ~ ( (22'h7ece <= (((2'h3 % (r90 + ( ( + ( 6'h1)) | $stime))) | r51) !== (27'h1d94 == (r189 & r252))))))) ? 2'h0 : r110))) <= ((r124 % r178) <= ( ( & ( $time)) - (((r22 == 27'h4da6) != 19'h14be) ^ (r155 / r52)))))));
		#10; r92 = (28'h4175 +  ( - ( ((( ( ~ ( (4'hf % (($stime ? 5'hf : ((((4'h8 | (r118 !== 10'h222)) != ($time / r53)) ?  ( ~ ( r49)) : ((r251 > r162) - r163)) == 17'h72a0)) && (16'h486b === r203))))) + r130) + 14'h3094) ? (((r153 | 12'h53b) + (((r97 ^ (28'h6257 > 4'h5)) !==  ( & ( ( ( ^ (  ( | (  ( & ( 13'h1537)))))) != ((18'h18c7 != r154) & r105))))) != r241)) - r193) : ((14'hcba !== (r26 | ($time && ((22'h643d ^ ( ( ~ ( r117)) < (r206 ===  ( ^ (  ( ! (  ( ! ( (11'h3b3 >= 27'h6d33)))))))))) / 6'h2c)))) > ((25'h6f8d >= 26'h4258) == ( ( & ( (( ( ! (  ( ~ ( ( ( | ( 32'h41ba)) + ( ( ! ( 14'h2b91)) + r190)))))) <= (26'h5532 + 14'h12cb)) == (r232 % ((21'h2891 / r76) +  ( + ( ( ( & ( ((8'h43 <= 24'h19c2) >  ( & ( 25'h70d2))))) + ((31'h65e0 !== (10'h18a ^ 1'h1)) < r191))))))))) / ((16'h16d0 ? 26'h5ce4 : (r66 ?  ( ! ( r127)) : ((((((18'h6d90 ^ 19'h2911) % (18'h5898 * 3'h0)) && $stime) !== ( ( & (  ( ~ ( 25'h56ef)))) -  ( | ( r124)))) *  ( | (  ( ! ( (r62 ? r238 : (22'h5c72 <= 28'h4c3))))))) !=  ( | ( 22'h388d))))) | (((( ( + ( r248)) !== ((r240 % 30'h5a83) - r4)) + 31'h131) || r147) & ((r36 | (((((15'h5184 > 29'h7846) + 15'h4959) ^ (r123 * r200)) / ($time &  ( + ( (8'hc8 & 9'h1db))))) > 5'hd)) / ((r86 > 29'h4da1) !== r118)))))))))));
		#10; r222 = (r106 * 32'h1826);
		#10; r88 = ( ( ! ( ((((r249 != 18'h6b91) >  ( ! ( ((r65 == r236) & 7'h59)))) ? r146 : ((r162 === $time) <= r135)) > (( ( + ( 32'h2513)) !== r252) || r147)))) <= ((32'h371b == r72) < 5'h1f));
		#10; r131 = r22;
		#10; r48 = ( ( & ( (((( ( - ( ((r9 - 30'h63a0) * r22))) |  ( - ( r212))) ^ 10'h1d5) ===  ( ^ ( 14'h2dbb))) % (9'h178 % (r241 !== ( ( | (  ( ~ ( (((21'h280 !== ((29'h1c0a - (1'h0 + 2'h3)) / (26'h2be2 * (r98 &&  ( & ( 22'hac0)))))) | (17'h5864 || r147)) <= (r51 ?  ( ^ ( r226)) : (r15 !=  ( | ( (8'hb6 && 6'h34)))))))))) < (9'h1bb != r114))))))) === r208);
		#10; r217 =  ( | ( (r7 || ((r98 === (r212 === ( ( ! ( $time)) | (6'h3 + 23'h6819)))) / (r154 >=  ( & ( r135)))))));
		#10; r145 = ((7'h5d > r79) !=  ( - ( r98)));
		#10; r22 =  ( ~ ( 22'h43eb));
		#10; r115 = r221;
		#10; r239 = (r198 !== (10'h79 !== (12'h444 ^ ((r204 && r214) %  ( ~ ( r7))))));
		#10; r170 = ((r185 % 25'h5b50) - r104);
		#10; r139 = (( ( ^ ( (((29'h158a && r170) ? r64 : 26'h4955) - (r100 >= r61)))) * r136) | r122);
		#10; r78 = 7'h10;
		#10; r72 = r70;
		#10; r145 =  ( | ( (8'h86 && r159)));
		#10; r123 = $stime;
		#10; r220 =  ( ! (  ( ~ ( ((((r79 === 12'hd3) && r55) % ((r1 <= ((r226 % (( ( | ( r107)) != r227) < (($stime < r242) !=  ( ! ( ( ( ! ( 29'h6b4e)) * (r221 || ( ( ! ( 29'h162a)) > 25'h45be)))))))) !== ((( ( ! (  ( | ( (r179 <= $stime))))) && 20'h7a52) & r249) < 29'h58eb))) & 25'h4a32)) == (r63 == r136))))));
		#10; r31 = 32'h3c62;
		#10; r216 = (r148 != r198);
		#10; r140 = r215;
		#10; r227 = ((r246 ? $stime : r163) && (((( ( ~ ( r157)) + 13'h1de6) / 2'h1) !== (($time <= (r195 &  ( ^ ( r121)))) && ( ( ~ ( r165)) * ((r124 !== 13'h9f1) && (r226 == (r79 <= ((r188 | ((((r70 >= (29'h4a7 % 2'h3)) < ((8'hba >= 4'h5) || 24'h394b)) !== r140) + $time)) / r68))))))) && r193));
		#10; r168 = 2'h3;
		#10; r208 = r211;
		#10; r196 = ((((r227 < 24'h299e) != 10'hac) && (((r16 && ((r10 ? ($time / $stime) : r229) >=  ( & ( (( ( | ( ( ( | ( 15'h5c9d)) /  ( ^ ( (r242 !== r117)))))) && r200) <=  ( & (  ( + (  ( ! ( r228))))))))))) - (7'h2c != (( ( & ( 17'hd65)) ^ $time) + (r82 >= r124)))) ?  ( ^ ( r222)) :  ( & (  ( ^ ( ((r146 != $stime) ^  ( ! ( (r4 %  ( ^ ( r114)))))))))))) ^ r88);
		#10; r200 = 12'h3e9;
		#10; r158 = (24'h2147 - 4'h4);
		#10; r72 = r219;
		#10; r101 =  ( | ( (r104 + r252)));
		#10; r98 = (27'h401a ^  ( | ( ( ( ~ ( 13'h74a)) * (( ( ^ ( r121)) ? 5'hf : ( ( ^ ( 17'h6a2d)) % 2'h3)) != (r43 === (32'h2ec9 %  ( - (  ( ~ ( (($time !== ((21'h583a +  ( & ( r117))) * r30)) <= r167))))))))))));
		#10; r57 =  ( ^ ( r87));
		#10; r54 = ( ( + ( ((( ( - ( r109)) ? 6'h9 : r99) - 28'h6c8c) + ((((((25'h46be && 14'h16f3) > r158) / r249) % (r168 || (r95 ===  ( + ( (((((r204 % $stime) <=  ( + ( (27'hb65 != 6'h1b)))) <= ((r139 && (11'h577 || 27'h5dbd)) + 1'h1)) || ((((13'h9d1 !== 22'h14cf) | (26'h101a + 23'h31a9)) | ((7'h4b - 26'h63f8) | (30'ha4d * 32'h760))) < ( ( ^ ( 3'h1)) < r111))) < (((r215 & 32'h4838) / ( ( ^ ( (24'h2d6f || 28'h4fde))) && ((4'hb <= 9'h24) & r112))) | (r97 === (r76 < 8'h76))))))))) ^  ( ^ ( ((26'h3743 || ( ( - (  ( ! ( ((3'h4 * ((7'h66 !== 32'h4200) & 14'h2b24)) ?  ( - ( r57)) : 21'h6ef))))) <= r70)) | ((r159 <= r181) - ( ( + ( (r36 || (r49 != (r185 ===  ( ^ (  ( ! ( 10'h2dc))))))))) === r150)))))) >=  ( | ( ( ( & (  ( ! ( 22'h416f)))) !== (r137 +  ( | ( $time)))))))))) ^ r148);
		#10; r44 = (11'h11 || 13'h99d);
		#10; r213 = r254;
		#10; r101 = 31'h6ed;
		#10; r190 =  ( ^ ( r133));
		#10; r222 = (32'h2008 >= 24'h68a3);
		#10; r12 = r13;
		#10; r235 =  ( + ( (r42 / $stime)));
		#10; r50 = ( ( ^ ( ((r251 <= ((27'h6eee >  ( & ( (($time ? r43 : $time) !== (7'h36 !== ((((((23'h6f4 != 26'h7c8b) & (32'h5eeb < 25'h6227)) | $stime) * (((29'h6a61 === 11'h6bf) & (30'h6956 / 21'h637d)) > r209)) +  ( | ( (($time % (22'h3516 ? 11'h405 : 6'h5)) % (11'h49d >= (4'he ^ 17'h9e1)))))) + r82)))))) & r152)) * ((((((r53 & r240) != ((((r146 === ((14'h1ccc - r221) % 1'h0)) !== ((( ( | ( 23'h24bd)) & r79) >= (26'h2a62 / 23'h59d6)) !== r94)) < ( ( ! (  ( ~ ( ((26'h1762 / 12'h3bb) ===  ( ~ ( 20'h2582))))))) > r104)) * r190)) != (21'h5a98 >= r53)) && ($time * 13'h1dc3)) / $time) - r217)))) < (( ( - (  ( + ( (2'h2 !== r32))))) != ( ( ~ (  ( & ( (r130 != ((29'hc97 - $time) ^  ( - ( r18)))))))) - r102)) + r33));
		#10; r224 = r199;
		#10; r74 = 31'he64;
		#10; r92 = ((( ( ^ ( ((r138 ? (((((r82 == (r128 * (r32 % (15'h7083 <= r219)))) >  ( + (  ( ~ ( 31'h75c7))))) && $time) <= 2'h3) | 23'h7c7b) : r20) + ((25'h4238 >= (( ( ~ ( r30)) < r97) ? (((((24'h5cda + r34) === 31'h60c9) != r72) == 11'h5c8) | (r92 / r77)) : (r26 != r174))) % (( ( + ( (((13'h507 + $time) < (r230 < r79)) / (( ( - (  ( & ( (21'h77de >= 21'h595c))))) & (6'h29 == r159)) == r120)))) ? (( ( ^ ( ($stime %  ( & ( (r44 ^ 19'h4868)))))) || 29'h425) != ((((((27'h3be5 <= 21'h73b3) >= 5'h1e) -  ( ! ( (24'h14b5 | 12'h81f)))) != (((31'h6c1a >= 7'h66) != (21'h2b37 * 5'hc)) | 26'h1e08)) ? $time : ((r238 && 9'he4) | $time)) / $time)) : ($stime || 10'h2af)) | 30'h6f3b))))) !=  ( & (  ( & ( (30'h2102 - (r214 ^ (r148 != r173)))))))) || r12) + $time);
		#10; r20 = (r109 ? (((((r205 * r142) - ($time && (14'h12d7 & (25'h300a ^ $stime)))) != 8'h46) ||  ( ~ ( ( ( + (  ( ~ ( ($stime <  ( ! (  ( ^ ( (r127 + r51)))))))))) == (r175 %  ( ! ( (((r70 == r189) > (((r1 !== 9'h40) != (5'h3 !== r198)) + (r221 ^ 30'h283b))) || 29'h1a0c)))))))) + (((r220 + (26'h5440 != (2'h1 == 6'h2e))) & r219) & 28'h5a06)) : (14'h1a0a < 6'h15));
		#10; r253 =  ( ! ( 32'h3419));
		#10; r95 = 16'h3cbd;
		#10; r49 = 2'h1;
		#10; r17 = (r251 <= r61);
		#10; r151 = 4'h7;
		#10; r136 = (r253 || ((r68 <= 30'h5ad3) != (3'h0 %  ( + ( 27'h5cc2)))));
		#10; r35 = (r153 & (r74 | ( ( & ( r94)) <= r72)));
		#10; r120 = (30'h3c55 + ((r48 || r173) & r231));
		#10; r214 = ( ( & ( (r168 % ((((28'h55b2 ^ ( ( ! ( 8'h4b)) === 11'h221)) < r217) != ( ( ~ ( ((r213 /  ( + ( ( ( | ( (((18'h5f95 * 8'h91) || (7'h17 & 16'h8ab)) && r127))) == 16'h5aae)))) *  ( + ( ((r109 == ((((18'h3972 + 25'h7165) == (4'h4 >= 7'h58)) * (6'h2a - (28'h4a9a + 16'h768d))) != (r130 !== ((11'h36b < 17'h7bb9) / 31'h65db)))) ?  ( | ( r139)) :  ( - ( 28'h5d29)))))))) !== (((15'h7581 < 5'hd) + ((((20'h61ac ^ r219) < 1'h0) | (r79 ^ r25)) * (r90 < $time))) -  ( ^ (  ( - ( (( ( + (  ( + ( r130)))) == (( ( ~ ( r200)) >= 24'h433) < 1'h1)) + 17'h7ce2)))))))) ^ (( ( & ( ((r161 +  ( & ( ( ( ^ ( r63)) * (((r201 & (13'h1fa9 || 2'h3)) *  ( ^ ( r103))) * r28))))) | 1'h1))) === $stime) >  ( ^ (  ( ! ( r165))))))))) >= ((( ( | ( 3'h6)) | r66) | 5'h8) ?  ( - ( r24)) : (r227 /  ( ^ ( ((( ( ~ ( (((r63 * ( ( & ( (r92 / (24'h565a + 12'h647)))) - (r124 < r138))) ||  ( - ( (18'h1d84 | ((r186 - 28'h4f76) | ( ( - ( 4'h5)) != 25'h57d1)))))) ^ ((r196 >=  ( | ( r186))) ? ((32'h15b6 & (26'h458a >  ( ! ( r103)))) / r171) : r99)))) || (($stime - (((((r64 | r129) / 18'h31eb) | $stime) & (1'h0 / r226)) !=  ( + ( r173)))) != r3)) % (r109 >= 9'h119)) + (((((20'hf4b ?  ( & ( (16'h394b > ($time *  ( + ( (16'h480 === 32'h42fb))))))) : 24'h56a7) ? 22'h5ab9 : r136) === 14'h2f0a) <= r83) % r134)))))));
		#10; r223 = (r227 ^  ( ! ( ((28'heb ?  ( + ( (r213 | (20'h18bc >= r78)))) :  ( & ( 10'h333))) | ((r132 != r21) - (r23 | r235))))));
		#10; r70 = $time;
		#10; r76 = (r49 / (((( ( - ( r188)) && r46) <= (r73 * r159)) || (r109 ^  ( & ( 13'h12a8)))) / (( ( - ( $stime)) > (r165 / ((25'h7b9e *  ( - (  ( ^ ( (((r28 + (r247 >  ( - ( (2'h0 % 10'h360))))) % 13'h48d) ? (29'h6a6f - 27'h5199) : 22'h2db7)))))) < 17'h6a8e))) >=  ( ^ (  ( - ( 5'h3)))))));
		#10; r184 =  ( & (  ( & ( r95))));
		#10; r244 =  ( | ( (12'hb7 / 9'hb9)));
		#10; r239 = 19'h7f7c;
		#10; r246 = (r224 != ((($time < 11'h493) !== (18'h148b - r178)) == (7'h4c < (r198 &&  ( | ( ((((((r140 &  ( ~ ( (( ( - ( 15'h988)) | r21) || ( ( ^ ( 11'h5c4)) <= (20'h7942 >= 15'hca5)))))) % r6) && (($stime + 6'h16) >  ( & ( 13'h76d)))) > ( ( - ( r13)) >= ( ( + ( 13'hc6a)) / (r247 * r180)))) >= (7'h20 || (( ( ! ( (((12'haae > 10'h15a) && 16'h4261) > r16))) & ((r100 / (r60 + (r99 / (27'h2093 - 8'hd5)))) - r234)) & ( ( ! ( $time)) === $stime)))) >= r31)))))));
		#10; r208 = r57;
		#10; r120 = 26'h5f9c;
		#10; r176 = 5'h2;
		#10; r205 =  ( ^ ( 31'h6209));
		#10; r219 = (1'h0 *  ( | ( r56)));
		#10; r9 = 19'h2d05;
		#10; r112 = ( ( ~ (  ( + (  ( ^ ( r163)))))) <=  ( - (  ( | ( (r78 % ( ( + (  ( ! ( $time)))) != (31'h4aff * r79))))))));
		#10; r163 = r143;
		#10; r20 = (((r127 | 17'h3217) ^ r11) || (8'ha2 != (r189 === r201)));
		#10; r45 = ((r171 ^  ( ! ( (r42 === 5'he)))) >= 13'h1b72);
		#10; r72 = ( ( | (  ( + ( r110)))) - 10'h189);
		#10; r238 = $stime;
		#10; r234 = r199;
		#10; r247 = r34;
		#10; r138 = r206;
		#10; r245 =  ( | ( r167));
		#10; r253 = (( ( | ( 14'h394d)) != (( ( ^ ( (((10'h1c6 == r212) ?  ( + (  ( ~ ( r148)))) : r51) ? ( ( ^ ( $time)) < r233) : (7'h3c ^  ( ^ ( 17'h7cde)))))) !== ( ( | ( r155)) !== r64)) <= r224)) % (( ( + ( (r79 === ((1'h1 <= (r81 / r68)) + (r139 != ((r180 ?  ( + (  ( ! (  ( ~ ( r46)))))) : (r171 % r237)) * r102)))))) %  ( ^ (  ( | ( r78))))) <= (17'h2b1f ^ ((17'h3160 ^ r59) > (((6'h3 + $time) * ((7'h3f !== $stime) ^ 3'h2)) ^ ((r181 > (r221 | (((r187 !=  ( - ( (((14'h3871 - 31'h1261) < (8'had / 6'ha)) & r192)))) || $time) ?  ( + ( r154)) : $stime))) +  ( & ( 21'hfbf))))))));
		#10; r193 =  ( & ( 15'h1a54));
		#10; r143 = r132;
		#10; r161 = ($time &  ( ~ ( (r107 ^ $stime))));
		#10; r47 = r197;
		#10; r72 = ((($time == 14'h3eb9) !== r242) < 12'hee0);
		#10; r167 = ( ( ! (  ( + ( r50)))) +  ( ^ ( (r231 * ((6'h26 <= ( ( ~ ( ( ( + (  ( - ( ((( ( + ( (2'h1 != 19'h3fa5))) === ((6'h11 % 4'h1) / (10'h37a / 30'h1e1c))) * 9'h1b6) != ( ( & ( (8'h22 === 2'h1))) * $stime)))))) * 13'h1daa))) * r192)) === 26'h5f03)))));
		#10; r99 =  ( ~ (  ( ~ ( r218))));
		#10; r66 = ( ( ~ ( ((( ( ^ ( ((11'h73f ? ($stime ===  ( ~ ( r187))) : ((((20'h4125 + $stime) | r85) == r13) === ((22'h47f0 & (r164 %  ( & (  ( + ( (23'h1879 + 19'h28f2))))))) >= 4'hf))) * $stime))) ===  ( ^ ( 29'h67cf))) ||  ( | ( r240))) >  ( - ( (r78 + (23'h272f && (r132 != (( ( & ( (($stime === (((16'hed3 * 1'h0) < $time) && ((6'h2 / 9'h101) ? (21'h637d - 26'h4190) : r63))) * ((((9'haf & 14'h2ce7) ? (2'h2 & 9'h197) : 9'hd5) <= ( ( + ( 27'h32c1)) && (9'h147 - 5'h11))) >= (r159 == (r200 <= 28'h3218)))))) ^  ( - (  ( + ( (r202 ? ( ( - ( 14'h190e)) % ((16'hffb >= 26'ha6d) + (23'h3a46 | 3'h4))) : r83)))))) % r246))))))))) ? ( ( ! (  ( ^ ( ((r117 === r65) & (r92 & r196)))))) / ((((((16'h4c37 !== ((r124 * r17) < (r161 + ((r55 === ( ( ~ ( r209)) & 10'h3fc)) % ( ( & ( ((7'h2f + 18'h274a) * (31'h4de5 < 12'hb26)))) >=  ( ^ ( ((14'h3161 >= 25'h7632) * (25'h2a76 * 8'he))))))))) >  ( ! ( ((10'h390 - r60) % (((13'h649 +  ( - ( r187))) !== r61) | 19'h40eb))))) >= (19'h49d9 <= r1)) & (( ( & ( r174)) == r111) / 18'h4732)) - ( ( ! (  ( | ( (r232 > r110))))) + (r73 < $stime))) <= r163)) :  ( ^ (  ( ! ( ((((r195 | ( ( | ( 22'h41f9)) ? (23'h754e / 6'h28) : (25'h7d32 == (4'h6 < 5'h1f)))) &  ( | ( ( ( ! ( r87)) - r71)))) -  ( ^ ( r179))) | ( ( & ( (3'h2 > $stime))) +  ( ! ( r165)))))))));
		#10; r9 = (26'h2a2e != 15'h83d);
		#10; r125 = 15'h6f76;
		#10; r245 =  ( | ( 28'h74c2));
		#10; r157 = r203;
		#10; r166 = ((21'h29d6 != (($time - r242) == ( ( & ( (((11'h323 &&  ( ~ ( (1'h1 + ((r68 / (((13'h18c8 + 15'h2554) % r147) === (9'h40 === (4'he || 1'h0)))) ^ ($time & r189)))))) | 30'h4919) <= r151))) < (r137 ? (r50 % (( ( - ( $time)) >= 19'hbdc) * r216)) : ( ( ~ ( (6'h3d | $stime))) <= 1'h0))))) <= ( ( - ( r229)) >= 22'h3540));
		#10; r138 = r246;
		#10; r163 = 32'h357d;
		#10; r251 =  ( & (  ( - ( r85))));
		#10; r83 = ((23'h34a0 <= r246) === 11'h66b);
		#10; r183 = (r152 || (($time ? (21'h6ca4 > 28'h650) : r140) != ($stime !== 27'h1214)));
		#10; r171 = 32'h6d44;
		#10; r180 = 9'h180;
		#10; r167 = (r199 ?  ( | ( r212)) : 23'h3844);
		#10; r221 = 12'h1b;
		#10; r198 = (r72 ?  ( ! ( r4)) :  ( - ( r213)));
		#10; r97 =  ( & ( 14'h290e));
		#10; r164 = 5'h3;
		#10; r33 = ((($stime || (7'h9 >= 9'h1bf)) < 14'hb12) < ((r246 / ((r116 ? 20'h1b7c : ((r189 + 17'h6013) - $time)) % $stime)) == (r100 ^ ( ( ~ ( (r189 !== r96))) & r40))));
		#10; r154 = ( ( - ( ((26'h562a && r20) && (r167 | ( ( & ( (r219 | (r185 ? (r114 || ($time / r206)) : (1'h0 < $stime))))) ^ 21'h4aae))))) /  ( ~ ( (r253 % ($stime * 15'h5c88)))));
		#10; r25 = (r5 & r139);
		#10; r205 = ( ( ! (  ( ! ( 29'h4196)))) && ((13'h19ed != (r149 != (24'h3ba0 !== ((r142 != (30'h3f71 || r189)) - ((((r109 / ((8'h1b % ( ( | ( r115)) ===  ( & (  ( | ( 30'h3325)))))) ||  ( + ( 6'h6)))) !== r180) || 26'h3874) - ((((15'h26a5 - ((((10'h36c % 18'h1c8) && (3'h0 <= 1'h0)) !==  ( & ( (30'h1ae9 - 29'h35cf)))) > 23'h24e9)) ||  ( & ( (r194 * r105)))) & $stime) %  ( ! ( (( ( + (  ( | ( r76)))) | ( ( ! ( ((3'h5 - 10'h2ec) + (32'h73bf & 20'h6da1)))) <= r79)) / r48))))))))) % r32));
		#10; r180 = ( ( | ( ((12'hc2a %  ( + ( (((4'he < r151) >=  ( ! ( r53))) >= (((( ( ! ( ((7'h1a ? ((21'h60e7 / 26'h652f) /  ( ! ( 16'h3871))) : (29'h69c9 && (29'h415d >= 15'h4e98))) && (((27'h4d27 === 5'h11) == (5'h7 / 27'h23f2)) >  ( + (  ( ~ ( 18'h3e82)))))))) != ( ( ! ( ( ( - ( r245)) != r141))) < (((r169 && 18'h2377) * ((19'hf5c && 21'h6ee0) || 2'h3)) / r178))) * ((((((16'h46dc >= 13'h54) >= (17'h793b >= 25'h35db)) < ((27'h7f99 > 23'h7718) != (12'hc9e == 3'h3))) || ( ( & ( (17'h2856 !== 18'h357))) * r241)) && ( ( ~ ( ((12'hfd6 * 14'h2446) / r102))) ||  ( ^ ( (r18 ? r25 : r123))))) == 5'h13)) ^ r185) | r245))))) !== (((r52 && ($time == r43)) !== ((14'h101e < ( ( + (  ( & ( ( ( + ( r195)) !== r50))))) ||  ( - ( 20'h140)))) != ((r48 != (r78 >= 6'h1c)) | (9'h8c ^  ( | ( 29'h4eb7)))))) < (((r199 + 11'h4f4) || r190) != 19'h5fcb))))) !== (((($time ==  ( + ( 4'hf))) /  ( + ( (24'h4ff8 * ( ( ! (  ( - ( (((((r11 | (11'h26b - 6'h39)) ^ r52) & (($stime % (15'h3778 == 15'h3a4a)) % $stime)) ?  ( ^ ( (r49 > r191))) :  ( ^ (  ( & ( ((15'h721d >= 11'h498) !== 13'h113c)))))) == r247))))) !== 15'h3ec5))))) === r154) |  ( & ( ((31'h5377 && ((r11 || ((((r70 > (r202 !== r43)) ? (r221 >= (((r255 == $stime) <  ( | (  ( - ( 23'h36a7))))) != (13'h1664 !== 32'h669a))) : r32) | (((7'h56 && 5'h1b) && (r106 == r168)) !==  ( & ( ((22'h15c7 && (r210 ^  ( - ( 30'h3a9c)))) ^ (((6'h12 | 1'h0) - (24'h3128 * 26'h265)) === (31'h947 | (28'h7be5 & 31'h336f)))))))) & ((r91 +  ( + ( 17'h1d47))) & (( ( | ( 28'h2f2)) &&  ( ^ ( 26'h663d))) <=  ( ~ (  ( ! (  ( ! ( (19'h5235 % (19'h3511 - 32'h5628)))))))))))) || (13'h82e | (r15 || (20'h145c != ( ( & ( r228)) == ( ( - ( (((2'h3 ? 10'h31f : 8'h32) +  ( & ( 13'h567))) % ( ( ^ ( 5'h2)) <= r117)))) != (r138 ==  ( & ( 14'h2b3a)))))))))) && (8'h99 ^  ( & ( (((((r157 + (30'h3c00 || $stime)) / r106) === ($stime !==  ( + ( ((9'h1b1 > ((19'h62e4 * 22'h2f20) - r190)) / 25'h38aa))))) != r200) % 1'h1)))))))));
		#10; r29 =  ( + ( 8'h46));
		#10; r70 = (r45 ? ((2'h0 >  ( & ( ((((28'h54b0 != ((r240 <= r248) - ((r123 <= 20'h4d70) ^ (r183 == (r182 ==  ( + (  ( + ( (11'h50f && 24'h6d05)))))))))) == (9'h45 %  ( & ( (20'h5daa | (((( ( + ( 7'h66)) && (23'h2117 && 5'h15)) ? r134 : 14'h2f50) > r236) != r231)))))) ? 8'hbc : ( ( ! ( (( ( | ( ((r70 * (18'h58fb ? r227 : (19'h4843 <= 23'h461d))) === ( ( + ( (7'h30 ? 13'h163e : 8'hb2))) & ((16'h7ef || 18'hef9) > (28'h3502 < 25'h15a7)))))) - 9'h1ad) - (((r129 | r81) > r41) || (r76 <= 17'h6b6e))))) &  ( | ( r125)))) <  ( + ( r6)))))) | ((r75 === (4'h3 !== (24'h4381 <= r157))) + r112)) : r244);
		#10; r146 = (( ( + ( ( ( - ( 16'h6078)) + (r112 -  ( | ( 26'h4c17)))))) <= (( ( - ( ((r203 | (((12'h954 ? ($stime |  ( ! (  ( - ( ($time && (9'h1b3 !== 19'h3078))))))) : $time) == 19'h4592) >= ( ( - ( $stime)) >  ( - ( 12'h242))))) >=  ( | ( ( ( & ( 32'h6a4c)) <= r3)))))) * (6'h14 ==  ( | ( r84)))) * (((((((11'h412 - r64) ===  ( | ( ((r141 ||  ( ^ ( ($time !== $time)))) ^  ( ~ ( $stime)))))) * r242) ? (31'h4adf | (r170 && (($stime * (r75 ^ (4'h3 < 23'h1faa))) >= 14'h2445))) :  ( + ( r186))) === r215) % r60) % ( ( & ( (4'h0 || $time))) ^ r179)))) > r82);
		#10; r219 =  ( | ( (9'h14b *  ( ^ ( ($stime ^ 12'h40c))))));
		#10; r164 =  ( + (  ( - ( 5'h18))));
		#10; r197 = (r243 % (( ( & ( r105)) && 25'h3a96) * (23'h1425 | $stime)));
		#10; r50 = (((r217 & r223) !== $time) + r81);
		#10; r185 = (5'h6 | (r31 >= r194));
		#10; r133 = (r210 / r112);
		#10; r203 = $stime;
		#10; r178 = (14'h258f <= 14'h1fb1);
		#10; r235 = ((12'h62a == ((r235 - r30) ^ 11'h49b)) ?  ( & ( 13'h1647)) : r237);
		#10; r46 = (r241 !== (((((13'h1466 ===  ( ~ ( (((r106 - r139) >=  ( ^ ( r97))) + 12'h69d)))) >=  ( & ( ((r94 ^ r251) <= 10'h389)))) && 28'h116b) <=  ( | ( ((( ( ! ( ((20'h14cc !=  ( & ( r45))) != r97))) + $time) == (( ( + (  ( ~ ( (11'h166 % (r79 ^ 15'h4c0a)))))) % ((27'h4742 + (r109 !==  ( ! ( (r238 >= ((13'h1bc2 ? 27'h21ab : 12'h85d) / r65)))))) ? (( ( - ( 22'h3a77)) && (r24 === (( ( + ( 24'h42f9)) <= (17'h1d1c >= 30'hed9)) -  ( - ( 31'h3f78))))) <= (r57 * (r252 !== r239))) : r117)) % r175)) === r66)))) ? ((r105 - r24) >=  ( & ( 6'h3f))) :  ( ~ ( ((((r27 || ((r72 != r105) === 30'h5332)) <= r58) < $time) > (r11 ^  ( & ( 28'h5de6))))))));
		#10; r14 = r60;
		#10; r158 = 3'h0;
		#10; r92 = 16'h5cb0;
		#10; r168 = (22'h238a == ((29'h737d % ((($stime || (r170 & ((((30'h2570 ? r246 : (r90 == (((2'h2 <= 11'hb6) > (20'h333a ? 3'h0 : 19'h4cae)) ? 8'he0 : ((16'h63a % 19'h22bd) - 12'h78c)))) != (r152 ? (r232 ? (((29'h7a19 >= 28'h28d5) ? (12'hdd9 + 19'h6d4d) : 16'h2ab9) ^ (r196 / (5'h6 >= 31'h55a4))) : r35) : r73)) <= (20'h4ff2 -  ( - (  ( + (  ( | ( 3'h0)))))))) % 5'h15))) * r34) !== $time)) ||  ( & ( 17'h1c43))));
		#10; r31 =  ( + ( ((3'h6 ^  ( ^ ( (r30 * r118)))) % ( ( - ( ((r131 <= r109) | ( ( - ( ($time %  ( ! ( 1'h1))))) + $time)))) / r228))));
		#10; r227 = r113;
		#10; r69 =  ( + (  ( | ( ((r175 * r252) >= 32'h458)))));
		#10; r160 = r171;
		#10; r99 = r171;
		#10; r26 = ($time >= (14'h3a77 ^ r235));
		#10; r188 = (( ( ! ( 19'hce0)) ^ (r32 ? (($stime <= (r90 * 15'h5bc5)) < r45) : (30'h7f25 == ( ( & ( ( ( ~ ( ((r137 / 22'h505) && r114))) || r72))) != r210)))) === (r220 | r130));
		#10; r210 = r221;
		#10; r241 = ( ( + ( r24)) + 10'h16e);
		#10; r24 =  ( + ( (3'h1 + 27'h6ef2)));
		#10; r104 =  ( + (  ( ~ ( r45))));
		#10; r39 = 12'h75f;
		#10; r136 =  ( - ( 5'h18));
		#10; r186 = $stime;
		#10; r202 = 3'h6;
		#10; r216 = 25'h70bd;
		#10; r208 = r211;
		#10; r143 =  ( + ( (r114 < r197)));
		#10; r118 = ((r187 * r55) <=  ( & (  ( - (  ( - ( ((( ( ~ ( 14'h3306)) % (((15'h67f + ($stime ^ ($stime %  ( ^ ( ((11'h82 < 18'h7222) ^  ( + ( 25'h1c3b)))))))) - (($stime <=  ( ! ( ( ( | ( (29'h166e % 7'h22))) >= 21'h608)))) <=  ( ^ ( ($time > r232))))) | r5)) > 2'h2) !== r89))))))));
		#10; r234 = 9'h1f5;
		#10; r254 = r6;
		#10; r39 =  ( & ( $stime));
		#10; r238 = ((15'h7bb7 >= 29'h70ec) & 22'hf47);
		#10; r65 = ((1'h1 - r123) + 12'h583);
		#10; r27 = (r221 == (r115 < r95));
		#10; r204 =  ( | ( 19'h10b));
		#10; r232 = (r78 /  ( ~ ( (((((8'hfa < r34) *  ( + ( (r91 != ($time + (3'h2 ? (21'h3c7a / r249) : (r205 * ((r71 % r26) && r39)))))))) | (1'h0 >= 21'h4545)) != 31'h1e16) !== (((5'hc / $time) == 27'h150d) !== 5'h1)))));
		#10; r213 = (r116 || ( ( ~ ( 9'h1cc)) !== (((23'h10fb == (((((21'h5703 * $time) >= ((29'h1274 !== ( ( - ( 11'h56d)) |  ( & (  ( + ( (6'h2 + 17'h129b))))))) >= ((( ( - ( r163)) > ((23'h2857 != 30'h64e4) / 5'h5)) || (((23'h7345 <= 21'hdf7) == r154) | r189)) > r117))) > (( ( + (  ( + ( r118)))) / 26'h7e4) <=  ( + (  ( - (  ( + ( (( ( ^ ( 16'h3752)) & (11'h2b && 4'he)) !=  ( & ( r63))))))))))) < ( ( ^ ( r82)) == ( ( ^ ( (( ( + ( $time)) ? ( ( ~ ( $stime)) > r142) : (13'h19ae | ((25'hced != 12'h2ff) !== 30'h290b))) && (r108 > r38)))) || (29'h7ef2 | r0)))) * $stime)) == ($time ? r49 : ((30'h1631 != (r225 - r55)) - (27'h3be0 ^ ($time ? 14'h2bb1 : r25))))) | 9'h1b9)));
		#10; r198 = ($stime <= ((2'h0 || (r230 * r145)) || ((r31 !== 20'h7fd3) !== (r98 %  ( ~ (  ( + ( (r110 <= $time)))))))));
		#10; r8 = 19'h16e0;
		#10; r145 = r147;
		#10; r125 = r193;
		#10; r182 = 1'h0;
		#10; r253 = ((10'h2de <= (25'h4a1d & r188)) < r181);
		#10; r44 = (24'h2e9a * (((( ( | ( ((r29 & r182) == r131))) / (15'h6295 | 3'h7)) > 14'had2) & r100) & (((7'h1b !== $time) % ((( ( - ( ( ( & (  ( + ( (r208 |  ( & (  ( + ( (1'h0 + 30'h6481)))))))))) / 10'h170))) != r170) === ((r216 && 20'h7e5a) || ((r115 &&  ( ~ (  ( & ( (r68 | (r149 < (r233 < r186)))))))) | r213))) || 15'h789)) && (r59 !== 8'hfc))));
		#10; r229 =  ( + ( r72));
		#10; r155 = 19'h69ae;
		#10; r56 = r65;
		#10; r84 = $stime;
		#10; r76 = $stime;
		#10; r235 = ((( ( ! ( r97)) | (29'h463 >= (( ( - ( r73)) | (r115 + $stime)) % 5'h15))) & ((r67 * ((( ( + (  ( ~ (  ( | ( (2'h0 !==  ( + ( (((6'h37 === 20'h7815) - (8'h25 & 26'h1ee9)) != 26'h152d)))))))))) % (r128 || (r140 *  ( - ( ((1'h0 > r41) == 17'h2448)))))) !== (12'h312 * ( ( ! ( r17)) > 6'h36))) + ((r172 ^ r139) /  ( & ( r127))))) || 29'h6f45)) ? (((r63 ^ ((($stime === 15'h3fb7) != (( ( ~ ( ((( ( ~ ( r77)) != ($time <=  ( | ( (19'h51cb != 19'hea0))))) ^  ( | ( (((27'h7fb1 ^ 22'h2e65) !== 8'h56) !== r60)))) + (8'h5b === (((10'h93 == r244) <= (14'h2620 && 3'h5)) <= ((22'h77e0 >= 13'hb60) &&  ( ^ (  ( ~ ( 20'h754a)))))))))) % ((((r106 & r242) | (9'h1a <= 17'h67c)) + ((r119 ^ (r206 < (r194 + (1'h1 <= 4'ha)))) ^  ( ~ ( r34)))) |  ( & ( $stime)))) +  ( ~ ( (r166 != 13'h147d))))) *  ( - ( ( ( ~ ( 3'h0)) %  ( ! ( r53))))))) ? (r102 == 3'h7) : (r60 * ( ( & ( ((r30 > (r33 <=  ( | ( $stime)))) ? ((r17 <= ( ( - ( 22'h7b0a)) ?  ( & ( (( ( - (  ( & ( 3'h0)))) & (r90 != (3'h1 !== 7'h2c))) / (((5'h14 ? 9'h1f : 21'h5421) & 27'h6fd6) ||  ( - ( r105)))))) : ((7'h52 + (r82 & (20'h218f !== (19'hca5 > 28'h7ddb)))) &&  ( | ( 15'h5da5))))) === 2'h1) : r187))) || 15'h3aa5))) & r178) : 16'h50d3);
		#10; r104 = r197;
		#10; r173 = 31'h818;
		#10; r205 = (((r254 >=  ( & ( (r51 || 10'h2bd)))) | ((12'h778 ? (4'h3 && ((r82 == r40) < ((r68 <=  ( ! ( ($time % r254)))) -  ( ^ (  ( - ( r179))))))) : (((r196 ^  ( ! (  ( + ( r61))))) == (18'h6246 < r0)) !==  ( | ( 23'h7fe)))) ^ r0)) & ( ( & (  ( | ( (10'h31a ? ((15'h5a76 != ((r49 > ( ( | ( (r106 % (( ( ~ ( 28'h4fd6)) -  ( + ( 29'h7066))) > ((27'hc41 === 28'hd4b) | (6'h2d & 8'h64)))))) && ((r242 <= 24'h2822) | $stime))) && r169)) != $stime) : r56))))) ^  ( | ( (r180 ^ r203)))));
		#10; r237 = (((((4'h5 -  ( ^ ( (((((((6'h27 ? ((2'h0 & 25'h3301) < (6'h25 | 9'h1ec)) : r223) | 31'h65e1) >= ((((31'h4659 + 17'h5965) <  ( | ( 11'h631))) !==  ( ~ ( $time))) * (($time / (10'h7d && 1'h1)) ^ 3'h1))) & 15'h5e87) ^ ( ( ^ ( r233)) &&  ( | ( 24'h3d10)))) == r49) >  ( - ( 2'h0)))))) - 5'h8) && 32'h3aa2) ? r27 : 27'h7c25) ? (25'h6fc1 !== (r8 & (((r82 >= 27'h5432) === ((25'h1d79 <  ( ^ ( 22'h53a7))) < r44)) / 2'h1))) : (r98 <= ((18'h56be === 13'h1971) % (r188 | r126))));
		#10; r72 = (r29 / ((4'ha - (( ( - ( ((r110 == (r68 != r28)) && 23'h1d5d))) !== $time) &  ( ! ( ((32'h122 >= r161) | 16'h36a9))))) < $stime));
		#10; r215 = r150;
		#10; r32 = (23'h22ba & r68);
		#10; r251 = ((((((((( ( & ( ((( ( + ( r230)) ||  ( ~ ( (10'h214 - 8'hca)))) & 29'h64fb) * r148))) <= $stime) == $time) - ((((((r247 >= r170) > ((r209 - r248) | ( ( - ( 15'h2d06)) ? 1'h1 : (14'h2f73 | 25'h3e87)))) % ( ( | ( r170)) > (r2 === ($stime > $time)))) !== r98) /  ( + (  ( | ( r156))))) +  ( + ( 30'h1f05)))) != r171) === (23'h16f4 & (((( ( + ( ( ( + ( ((10'h176 % 27'h709d) !== r155))) ||  ( ^ ( ( ( & ( 8'hbc)) !=  ( ^ ( 18'h426a)))))))) === r80) !== 23'h72f3) != r118) ^ (r122 -  ( ! ( (r57 * (25'h14f1 === (r168 / r149))))))))) | (r65 / $time)) == r250) ? r193 : r163) && 32'h1880);
		#10; r16 =  ( - (  ( - (  ( - ( r182))))));
		#10; r82 = r63;
		#10; r173 = 30'h254b;
		#10; r120 = (14'hd78 ^ r193);
		#10; r133 = ((r37 != r131) ^ r221);
		#10; r215 = ((25'hb1f || ( ( & ( (((((r198 | ((28'h6191 / 4'h2) >  ( & ( ((((25'h4f79 | 26'h5a16) ^ (3'h2 > 21'h51e3)) * 21'h31e8) >= (r25 / 26'h3a40)))))) !== (r33 %  ( - ( (((((15'h2a8c % 1'h0) + 32'h5653) + r172) || $time) ^ 23'h5215))))) == r173) != (23'h1aaa == (13'hccb ? r24 : (r86 && ((( ( ! ( (r126 !== (28'h2588 == 29'h7d09)))) == (24'h10c2 > 22'h5f23)) ||  ( ! (  ( - ( r16))))) % ( ( & ( r0)) ^ r129)))))) <= 3'h0))) - r115)) &&  ( ^ (  ( + (  ( ^ ( $stime)))))));
		#10; r98 = r156;
		#10; r129 = (((r44 <= (((r14 >  ( - ( r236))) < ((23'h5704 > (r163 === ((r136 != ( ( | ( 16'h7a29)) >= 21'h19b8)) !== (31'h53bd <= r38)))) !=  ( & ( 24'h332a)))) > (((((((r75 >= 23'h659f) !== (29'h2824 > r29)) <=  ( + ( r103))) - (r69 * ((r222 !=  ( & ( r11))) <= $time))) || (r252 - r29)) >= (9'h0 != 30'h7bb1)) ||  ( ^ ( (r204 != r33)))))) + $time) & (( ( ~ ( r161)) == 18'h371b) - ( ( + (  ( + (  ( + ( ($stime > 10'h349))))))) == $time)));
		#10; r224 = (25'h3bb6 ^ ((r169 !==  ( + ( (($time <= r231) ? 12'h7e7 : ( ( ^ (  ( ~ ( r186)))) >=  ( ~ ( ((r202 &&  ( & ( (11'h3f4 > (r148 < 24'h6a71))))) <= r104)))))))) == (((2'h2 % (((r226 < 2'h3) | (((2'h0 + (8'h1 || 7'h52)) !== ((r234 | ((( ( ! ( 12'h2fa)) + 23'h54ed) >=  ( ! (  ( - ( 6'h1e))))) >= r230)) != 20'h7209)) - (14'hc55 % (r243 != r235)))) & (10'h110 > r103))) ==  ( ! ( r102))) || $time)));
		#10; r15 = r135;
		#10; r18 = r148;
		#10; r179 = 13'h807;
		#10; r144 = r116;
		#10; r100 = r116;
		#10; r44 = $time;
		#10; r133 = 8'h67;
		#10; r119 = $time;
		#10; r155 =  ( ! (  ( + ( r55))));
		#10; r241 = (r252 == ($time || r154));
		#10; r162 = 21'h4542;
		#10; r154 = 25'h3c0a;
		#10; r172 =  ( & ( r130));
		#10; r152 =  ( ~ ( r25));
		#10; r229 = r1;
		#10; r238 = $stime;
		#10; r180 = 21'h942;
		#10; r231 = r199;
		#10; r39 = r247;
		#10; r46 = (23'h5bc != 3'h0);
		#10; r166 =  ( | (  ( | ( (13'h8cd ^ (((r12 || ( ( | ( 10'h14b)) && 12'h430)) === r195) & (30'h28c0 %  ( ~ ( 27'h521b)))))))));
		#10; r23 = r20;
		#10; r102 = ( ( | ( r216)) | 27'h7337);
		#10; r223 = ((1'h0 > $time) % r228);
		#10; r42 =  ( ^ ( ((r181 === r129) && ((r204 !== ((r112 ^ ( ( | ( 9'h199)) <= (r75 == ( ( ! ( 28'h5b63)) <  ( ~ ( ((r96 <= (((15'h6ad0 !== 13'h5a1) <=  ( ~ ( 24'h2def))) == ( ( ^ ( 24'h146e)) / (28'h13b1 >= 11'h94)))) ||  ( + ( (( ( ! ( 27'h51f3)) >  ( & ( 10'h2c7))) -  ( ^ (  ( ! ( 1'h0)))))))))))))) == ( ( ^ ( (( ( ^ ( (((32'h4dc3 - (r216 - 27'h503c)) <= 11'h1fd) |  ( | ( r46))))) && 22'h5f72) === r74))) !== (r190 / ((r33 ||  ( | ( ( ( + ( r53)) !== (28'h1cb9 || ( ( | ( (1'h1 && 27'h699))) *  ( & ( (16'h3dd0 === 17'h5fae))))))))) ^  ( | ( 12'h1de))))))) < r38))));
		#10; r174 =  ( & ( 12'h666));
		#10; r79 = ((r135 && r189) !=  ( | ( r186)));
		#10; r150 = (3'h3 * ((r251 !== ((9'h1ef - $stime) - (( ( - (  ( - ( r49)))) || r241) == ((( ( - ( 32'h4db1)) == ((r247 !== ((($stime + ((16'h42ad != 23'h2b27) ? r203 : (17'h2b91 % 27'h7fd3))) + ( ( & (  ( | ( 12'ha1b)))) !== ((21'h4286 % 22'h536e) ^ 16'h6608))) ? $stime : 14'h380a)) |  ( ~ ( ((r115 & ((r16 + (30'h5605 & 17'h245)) - 19'h4ee4)) !== 14'h899))))) != ( ( ! ( r204)) >= (r58 + ((1'h0 === 8'h8b) + ((((9'h10 === r7) / r217) <= 5'ha) * r254))))) == ( ( & ( 6'hd)) && 11'h440))))) ^  ( - ( (r27 & ((r177 === (r226 != $stime)) | 9'hf))))));
		#10; r248 = r209;
		#10; r5 = r51;
		#10; r21 = 12'h97c;
		#10; r51 = ( ( | (  ( ! ( (r174 > ( ( - ( 8'h2a)) >= ( ( + ( (( ( ~ ( r65)) + 8'h41) ^ 28'h7bc3))) / (13'hf60 * r126)))))))) >= ( ( - ( $stime)) <= ((r14 ^ (r25 >= 10'h344)) & ( ( - ( 21'h2549)) <= ((22'h7049 > 4'hd) ^ r172)))));
		#10; r158 = (r89 !== (( ( ^ ( ((r215 <= r205) * ((r142 % 15'hce6) < r253)))) | r84) +  ( & ( (r75 >  ( - ( ( ( ! (  ( | ( (r183 > 26'h7d82))))) >=  ( ~ ( (((r79 % ((r124 === ((r168 *  ( ~ ( 19'h6332))) <=  ( + (  ( + ( 32'h4365)))))) & ( ( ! (  ( - (  ( + ( 31'h67f5)))))) && r70))) >= (1'h1 & ( ( | (  ( ! ( $time)))) !=  ( & ( 7'h57))))) + r71)))))))))));
		#10; r180 = ((r27 ? ($time -  ( - (  ( ^ ( r86))))) : r20) - (( ( ~ ( (( ( ~ ( (30'h1d1e == ($time == (23'h196b === r86))))) & (21'h7750 >= ( ( ~ ( ( ( ! ( ($stime == 25'h47c6))) % ($stime && r93)))) / ($stime && ((r237 || r84) ^  ( | (  ( + ( r121))))))))) %  ( - ( ( ( + ( r158)) + r54)))))) == ( ( | ( 16'h315f)) >= ((((( ( + (  ( ~ ( r74)))) + 20'h7b7f) ||  ( & (  ( + ( 23'h4708))))) | (( ( & ( (4'h6 === r209))) || 13'h9c8) / r229)) ^  ( | ( ((4'hf ? 24'h4865 : 16'h6051) > (10'h250 <= 16'h354))))) || (r139 === (6'h3e <= 16'h59a))))) || (r80 ? (($time !=  ( ~ (  ( ~ ( (r243 ? ((28'h741c % r164) +  ( & ( ((( ( & ( r252)) || 26'h14dd) && r76) % r123)))) : 12'h35b)))))) ? (18'h36a6 === r202) : (((((27'h473b | r219) * r121) | (r30 >= (( ( ! ( 21'h52b8)) != (3'h0 <= (r38 % (((4'hf === 17'h45ca) %  ( - ( 15'haa3))) === ((20'h6ddf > 31'h6ad1) !== $stime))))) < r48))) > r110) >= 6'h3d)) : r163)));
		#10; r72 = (( ( ~ ( ( ( ~ ( ( ( - (  ( & (  ( ^ ( r217)))))) | (r180 == r234)))) <= 24'h480a))) % $stime) !== (24'h5c74 > ((r244 | ( ( ~ ( (((((23'h971 /  ( | ( (13'h121f <= ( ( - ( 28'h6b51)) >= (12'hcfc || 2'h1)))))) ? ((r11 |  ( - ( 32'h450d))) > r254) :  ( ~ ( $stime))) + (r74 & r104)) ||  ( - ( r235))) | ((12'hafb % r158) - 17'h7d6b)))) ^ r225)) ?  ( ! (  ( ~ ( ((((((((((29'h532 <= 16'h3d4b) ? r138 : r213) || (16'h52cf > (10'hc9 + 1'h1))) || $time) >= 16'h2a91) |  ( & (  ( ^ ( r43))))) <  ( ^ (  ( | ( (r91 | 2'h3)))))) / r186) * ($time / (r182 != r171))) < (( ( ! ( 19'hf53)) % r173) ^ r90)))))) : $stime)));
		#10; r162 = (13'h1684 !== 20'h5bae);
		#10; r125 = $time;
		#10; r65 = ((21'h5040 %  ( & ( (r168 / (r250 * r214))))) <= (21'h5bf !=  ( ~ ( $time))));
		#10; r132 = 14'h1f62;
		#10; r35 =  ( ! (  ( - ( (((((((8'h0 % ((( ( - ( ((17'h4f6 || 23'h241d) * (24'h3ec2 <= 31'h7ec8)))) / $time) >= (r114 & r213)) == (10'h33f === r79))) ?  ( ~ ( 16'h7540)) : ($stime || ((r144 - 20'h7607) !==  ( & ( 6'h7))))) == ( ( ~ (  ( ^ ( (r251 / ( ( ~ ( $stime)) < (((12'hcdd & 7'h6f) && (18'h7be < 16'h51a7)) || ( ( ! ( 31'h5b74)) ^ r127)))))))) + r254)) - r158) ===  ( | ( 11'h317))) ^ (r88 -  ( ^ ( (( ( ^ ( r179)) | ((r137 <= r77) === ($stime == ( ( + ( (r190 !==  ( ! ( 24'h667d))))) ^ $time)))) / r135))))) | (((r151 ||  ( ^ ( $stime))) >= r38) == (((( ( + ( ( ( - ( 3'h5)) > (((((11'h7ed > 23'h4848) + (12'hbf8 / 5'hb)) ^ r115) && ((32'h4a9d | (30'h66c5 & 30'h3e62)) >= 22'h14fe)) > (((r54 | (19'h3af4 ? 20'h63c8 : 3'h6)) | ((5'h19 | 2'h0) >=  ( ~ ( 2'h2)))) === ( ( ^ (  ( ~ ( 5'h1d)))) != (r8 == (27'h69be % 32'h3b05)))))))) > 17'h6896) <= $time) * 9'h17e) >= (r253 | r11))))))));
		#10; r42 = 16'hf15;
		#10; r139 = ((( ( & ( (14'h3f9d ===  ( ^ ( 21'h5f2f))))) + 2'h2) % 22'h5b3c) !==  ( | ( ((( ( ! ( r51)) / r88) ? 9'h1a3 : $stime) > 9'h194))));
		#10; r8 = ( ( & ( 20'h40b8)) ? ( ( + ( (( ( + ( ($time | ((3'h4 <= r197) == r234)))) != r4) - (r114 * 23'h46dc)))) % r68) : r172);
		#10; r181 =  ( - ( ($stime % (23'h1d8f &&  ( - ( ( ( ^ ( $time)) | (r108 & r26))))))));
		#10; r159 = (((18'h535a % r30) * r65) >= ((( ( & ( ((((((r105 || 31'h4634) * ((r174 == (r61 ||  ( & (  ( + ( 6'he)))))) <= r233)) / $stime) || (((20'h55e8 * 20'h57da) != 27'h10ab) && (((( ( ^ ( (25'h574b != 25'h59bb))) % ((5'h13 === 17'h4256) !== (28'h5ecc !== 1'h1))) <=  ( | ( r173))) !== $stime) || (( ( ! ( ($time >= (12'h42c | 23'h60eb)))) % (($stime >= 14'h23de) == r219)) > r65)))) && (18'h7c43 !== r96)) != (( ( - ( ( ( - ( ((r100 ?  ( & ( r142)) :  ( - ( r30))) === r236))) <  ( ! ( r38))))) | $stime) - (( ( | ( r68)) <  ( ^ ( (29'h6ea5 === ((((10'h243 === 31'h625f) >  ( ~ ( 26'h75a))) - r95) <=  ( | ( (r92 === $stime)))))))) >  ( & ( ($stime >= r76)))))))) | r92) ^ (10'h2f2 !== $stime)) >= r103));
		#10; r35 = (31'h1e3a * 13'h289);
		#10; r50 = ( ( + ( ( ( - ( 13'h1945)) &  ( | (  ( ! ( r128))))))) * (((($stime >= 7'h61) || (((( ( ! ( (r180 > r44))) * (($stime >= (( ( + ( r106)) ==  ( ~ ( 32'h59e7))) || 5'h9)) && 13'hcd)) < ( ( & ( 15'h5791)) ===  ( + ( ($time - (((( ( ~ ( 30'h6092)) & r184) + 31'h27e1) == ((31'h1dfa + 7'h68) !=  ( ~ ( 22'h10ab)))) & (16'h30ab / r158))))))) ? 12'hcb7 : (31'h4c6d !== (26'h4e33 < ((20'h1dcd / ((( ( & ( (23'h3c7c < 4'h6))) % ( ( | ( 18'h6b37)) / (31'h56e7 - 9'h1b5))) - r174) >= 12'h281)) !== (r100 * r11))))) ^ r201)) *  ( | ( 21'h41a0))) <= r130));
		#10; r17 =  ( & (  ( + ( r76))));
		#10; r99 =  ( ~ ( ((((r50 + (((r49 / (($stime * $stime) >=  ( | ( r137)))) > (r27 <= 9'h151)) / ((((((r222 > r101) % r93) +  ( ^ ( (3'h2 ||  ( - ( 28'h2340)))))) == ( ( ^ ( (r62 | (r201 === $time)))) <= 18'h6c9e)) >  ( | ( r235))) <= ( ( ^ ( (((22'h402 | 12'h9b) | r92) * (r181 / ((r17 & $time) > r160))))) != r20)))) & (((r109 >= ((r237 == ( ( + ( ((((27'h7c62 > 5'h10) || 28'h4e87) | ((17'h62af === 21'h4f4) <  ( ! ( 22'h4838)))) >= $stime))) && 23'h2eb3)) ^ ( ( ^ ( (r112 < (r212 > 6'h3d)))) ^ ((( ( + ( 8'hcc)) && 22'h6bf5) >= (r109 <= (((8'h3a == 25'h11d) == 19'h19b8) /  ( & ( $time))))) ^ (32'h174d % 31'h75c7))))) / ((r37 >= ( ( ! (  ( ~ ( (r0 <= ((r215 * 27'h649a) + 20'h7c51)))))) < r221)) !==  ( ^ ( r159)))) === r133)) + (23'h38d1 ? ((($stime ?  ( - (  ( - ( ( ( & ( ($time < r66))) ? r170 : (( ( ^ ( ((20'h6ff5 * 26'h4341) - r78))) / r196) < r246)))))) : ( ( + ( ( ( | (  ( ^ ( 18'h3e9)))) ? r129 : r245))) %  ( ! ( r128)))) / $time) * r156) : 16'h1426)) == 9'h114)));
		#10; r102 =  ( ^ (  ( ^ ( ((r211 ^ (r229 === r249)) < (((r17 * r174) * r229) <= ( ( & ( 26'h56cf)) || $time)))))));
		#10; r7 = r109;
		#10; r195 = (r100 - r246);
		#10; r248 =  ( ! ( ((r14 === (((r120 > ( ( | ( r100)) !==  ( ! ( 2'h2)))) > (( ( & ( 6'h18)) %  ( | ( 1'h0))) &&  ( + ( r251)))) /  ( ~ ( ((r233 - 24'h7a6a) / r56))))) === ( ( - ( r104)) !=  ( ^ ( 1'h0))))));
		#10; r160 = r14;
		#10; r164 = r57;
		#10; r26 =  ( ~ ( r63));
		#10; r20 = 27'h7948;
		#10; r33 = (((r235 > ( ( + ( ((22'h4078 % 28'h43d5) ^ ( ( | (  ( + ( r216)))) == r196)))) || (((14'h3a11 - $stime) == ((r45 - 5'h5) ^  ( ~ ( ( ( + ( (((((11'h70b | 19'h604f) > (29'h2b8 * 4'h8)) ^ r130) && ( ( & ( (13'h2b5 - 14'h34f9))) ^ ($stime < 10'ha5))) < r19))) * (((( ( ^ ( (7'h51 === 9'h7d))) /  ( & ( r242))) *  ( + ( (r120 * (31'h3f97 != 27'h5c58))))) & 6'h2f) < ( ( & ( r148)) ^  ( + ( 14'hfd5))))))))) ==  ( ! ( r231))))) + r248) && ((r48 | (r187 | (r221 == ((r42 & r204) == r140)))) < r15));
		#10; r221 = (16'h49d1 || (r58 + ( ( + (  ( ^ ( r240)))) > r5)));
		#10; r245 = ($time | $time);
		#10; r80 = r72;
		#10; r47 = $stime;
		#10; r43 = r104;
		#10; r128 = r105;
		#10; r253 = r67;
		#10; r145 = r81;
		#10; r126 = 15'h9eb;
		#10; r24 = r162;
		#10; r233 = $time;
		#10; r182 =  ( ! ( (($time ^ (r171 === 11'h452)) - r95)));
		#10; r94 = r219;
		#10; r231 = (((((r234 == r75) -  ( ^ ( $time))) | ( ( & ( ((((( ( + ( ((((19'h3cbc != 29'h50b3) === r179) === $time) >= 31'h7c7b))) > ( ( & ( ((r174 & (3'h0 - 18'h4c8f)) / 23'h16fc))) !==  ( | (  ( ^ ( ((32'h1b5c * 24'h1c03) > r120))))))) || (( ( ^ ( r53)) != ((((8'hec <= 9'h169) !== $stime) === ( ( - ( 16'h304e)) < (26'h3834 <= 18'h58bc))) ? 25'h6ca3 : 27'h60a2)) >= 7'h74)) - $stime) !== ( ( & ( (r193 <= r106))) &&  ( & ( ((9'hc || r173) != r85))))) /  ( ~ ( ((r82 / 25'h5809) <= ((r166 % (10'he3 -  ( ! ( ( ( ~ (  ( + ( 21'h5ea1)))) ? 32'h6caa : $stime))))) === (($time !== 15'h2f0c) > ((r134 && r13) & r131))))))))) < ((19'h706d && ($time & (($time === 18'h786a) <= 13'h1ed6))) ? (r176 == r217) : (r15 < (19'h4b23 ^ 20'h3584))))) ? 19'h46f1 : 16'h10bc) ^ (28'h57a5 >=  ( | ( $stime))));
		#10; r64 = (((( ( & ( ((((19'h1c36 >= 27'h1fc7) ^ r191) <= 18'h479f) && ((((((17'h38f5 / 16'h7871) > r19) <  ( ^ ( ( ( ! ( r255)) <= ((r196 / $time) ?  ( & ( r91)) : $stime))))) - (15'hc67 ^ ( ( ! ( (( ( | ( 10'h2bd)) == (9'hba > 4'h8)) + r104))) >=  ( & ( r46))))) !== ( ( & ( r158)) - (( ( & ( 27'h5bca)) ^  ( ~ ( r185))) === (r208 |  ( ! ( (((31'h3393 && 24'h16f4) <= (14'he7a / 15'h3c50)) & r73))))))) != ( ( ! ( 5'h14)) >= ( ( ^ ( 25'h2f7f)) / r25)))))) + ((7'h32 ^ (( ( + ( ((((r171 ==  ( - ( (24'h24c9 != 27'h188c)))) % (21'h1cd3 !== ((21'h4f82 !== 5'h5) !== (30'h592c && 31'h4d6)))) & ( ( | ( 32'h10e6)) * (r51 < (2'h3 &&  ( ! ( 9'hb5)))))) >= ((( ( - ( r100)) + (r94 < (4'h9 - 19'h7687))) / 30'h3d99) < ((22'h1717 <= (30'h7a58 ? 23'h26de : (2'h3 * 32'h15f2))) + r226))))) || r220) ^ r147)) & r163)) && 25'h4a4b) === r71) | 13'h13da);
		#10; r247 = ((r64 >= (6'h6 - 30'h1466)) < 10'h89);
		#10; r80 = 19'h4198;
		#10; r186 = r249;
		#10; r95 = r153;
		#10; r32 = 17'h76a7;
		#10; r81 = ((r230 & r127) >= ( ( ^ ( r166)) == (20'h625d % r106)));
		#10; r150 = r47;
		#10; r16 = ( ( ! (  ( - ( r127)))) == (20'h2d74 ^ ((( ( & (  ( + ( ($time ===  ( | ( r121))))))) - r238) | ((26'h7f81 | r147) || (16'h564f & r121))) | 29'h30a3)));
		#10; r159 = 7'h5;
		#10; r50 = r178;
		#10; r198 = (( ( ! ( $stime)) <= 30'h3341) >=  ( ~ ( (14'h2cc8 && ((((r238 ===  ( - ( ((18'h3731 || (21'h6044 > r225)) + $stime)))) && $stime) < ( ( - (  ( & ( ( ( + (  ( ~ ( 31'h5c4f)))) * r224))))) / (( ( | ( 17'h3bc0)) / r141) & r154))) ^ ((r176 + ((18'h3d71 === r214) ^ ((($stime >= r179) |  ( + ( 6'h28))) % ((r91 + ((r10 <= ($stime %  ( ! ( $stime)))) & (( ( & ( (24'h274b + 5'h1e))) == 30'h4efa) - (r23 > r185)))) !== (((r236 <=  ( ~ ( ($time ? (20'h6978 > 25'he4c) : (29'h18de | 13'h19a7))))) & (($time > ((27'h7cd5 || 10'h2d1) /  ( | ( 7'h69)))) != (((18'h6172 | 19'h59d4) == (30'h4c9b && 19'h2001)) !== ((15'h73ea % 20'h1953) ? r244 : r76)))) % (r143 ? (r59 >  ( ^ ( r141))) : ((19'h13f7 <  ( ^ ( (26'h7eda ^ 1'h1)))) != r136))))))) && $stime))))));
		#10; r100 = (((($stime ? r212 : ((r115 >= 13'hd24) === (( ( & (  ( + ( (( ( + ( r7)) != ((((17'h3105 ^ 16'h5f7b) != 28'h7cd2) && 7'h2) / ((r122 ? (20'h5bb0 != 26'h66d1) : (32'h251d * 30'h1913)) === r221))) / 4'h6))))) ? ((r54 && (24'h50eb / 3'h0)) - (r249 | r87)) : (( ( ^ ( ( ( ~ (  ( - ( ((18'h165 !== 18'h7eb7) || (29'h26d4 && 5'h6)))))) && (r36 <= (r140 % ((13'h1b93 && 10'h97) - (9'he6 % 10'h30e))))))) *  ( ! ( ((((4'h3 && (14'h151b || 32'h7a7e)) * r208) %  ( ^ ( r215))) <  ( ^ ( 29'h2bb1)))))) + ((r123 <= 29'h381e) >= ((r177 <= $time) && 22'h6707)))) > r183))) <= (((30'h2485 > (7'h5b * (((r8 != 27'h4ad2) & r75) == r104))) & ((r222 + r255) + 2'h1)) > 7'h48)) < r195) & (r232 +  ( - (  ( | ( 5'hc))))));
		#10; r111 = $time;
		#10; r220 = ( ( & ( 32'h47c4)) != ( ( ~ ( (($stime <= $stime) >= (r22 !== ( ( | ( 15'h82b)) | r125))))) - 20'h65a5));
		#10; r103 = ((r212 & (r10 != (2'h2 | (r201 -  ( ! (  ( ^ ( (r100 && (r69 % (r86 + 25'h2418))))))))))) % ((5'h5 || 3'h7) & (( ( + (  ( & ( (r236 + ((r25 &  ( & ( ( ( ~ ( (29'h682e +  ( ~ ( (23'h4ffa % 5'h7)))))) == 32'h6eb2)))) < r202)))))) ==  ( ^ ( 7'h56))) % (32'h14d5 +  ( - ( ((3'h7 | ((((( ( - ( 27'h237d)) !=  ( | (  ( | ( 25'h1e5a))))) ^ ( ( ^ ( (r244 === (28'h502d - 32'h2e48)))) / (r147 < r167))) && r42) > (( ( ^ ( (((18'h3679 === 24'h3b03) * (1'h1 - 17'h6b4)) | 3'h1))) != r141) < ( ( + ( 30'h1484)) &  ( | ( (((6'h3b === 20'h4cb9) % (23'h7809 !== 5'h7)) > 23'h79ca)))))) <= ( ( ! ( r254)) - r79))) <= ( ( + ( (r25 && $time))) % ((((22'h51e6 && (r206 * $stime)) !== r38) | r148) - r127)))))))));
		#10; r55 = r221;
		#10; r206 = r156;
		#10; r180 =  ( ~ ( 16'h2225));
		#10; r67 =  ( + ( (((r203 && r69) === r123) != r202)));
		#10; r75 = (( ( | ( ( ( | ( r9)) < (11'h3d9 ===  ( ! ( ( ( ^ ( r99)) === r224))))))) == 28'h2fb6) && ((30'h8c3 - r134) < 23'h5849));
		#10; r217 = (18'h2761 % (r56 | (($time < (20'h6ce0 *  ( - ( (r235 * (( ( - (  ( | ( ((((6'h3a + 29'h3b2e) == 12'h6d5) + r79) > (r156 && ((26'h257f == 2'h2) || (9'h72 == 16'h41d9)))))))) * ( ( ! ( ((r48 -  ( + ( (2'h3 + 14'hb38)))) ? r166 : r136))) !==  ( | (  ( + ( r74)))))) != ($stime > ((26'h39cb !== r112) % ( ( - ( r124)) == r221))))))))) < r23)));
		#10; r14 = (r167 <=  ( ! ( (r106 >= r22))));
		#10; r254 = (r246 + ((((r132 && ((( ( + ( 6'h0)) < r228) === (25'h5358 === ($stime % 15'h7d8d))) == r28)) || $stime) ^ (r24 *  ( ^ ( 13'h402)))) && ( ( | ( ((r100 + $time) === r249))) != ((19'h52e8 - 16'ha15) & (((1'h0 <= 23'h39c8) % ((19'h3f6b > ($time & r181)) >= r47)) + (( ( + (  ( | ( 2'h2)))) === r63) == r48))))));
		#10; r231 = $stime;
		#10; r198 = ((13'he17 === (( ( ~ (  ( ^ ( (r249 ===  ( | ( ((( ( ~ (  ( | ( ( ( ! ( 24'h53e3)) & (21'h3e5d != 22'h7f09)))))) >= r72) == r147) >  ( & (  ( ~ ( (7'h5c == r217))))))))))))) != r206) && ( ( - (  ( & ( (r203 / r196))))) & ($stime ^ ((7'hf && 6'h13) < 31'h2e8e))))) <= ((r29 >= r103) == 29'h4b73));
		#10; r208 = (r245 * 21'h176);
		#10; r232 =  ( ! (  ( ^ ( (r195 <= r240)))));
		#10; r120 = $stime;
		#10; r25 = $stime;
		#10; r36 = (( ( | (  ( - ( ( ( | ( r63)) & (( ( | ( 10'h279)) % ($stime != r51)) != ((( ( ! ( r108)) ? (r28 && (r75 / 13'h302)) :  ( | ( (r19 == 27'h2750)))) - (r135 + r97)) || $stime))))))) &&  ( & ( 29'h78e2))) >= 9'h9c);
		#10; r126 = 27'h5db1;
		#10; r7 = 27'h61d3;
		#10; r254 =  ( ^ ( 6'h32));
		#10; r76 = r9;
		#10; r106 = r11;
		#10; r115 = ((r69 > r37) && (r35 == r169));
		#10; r190 = r31;
		#10; r39 =  ( + ( (15'h2c29 ? r216 : ((13'h928 != ((r216 | r94) /  ( ! ( (r8 !== (r209 & 8'hc6)))))) + 29'h1e5d))));
		#10; r77 = r166;
		#10; r211 = r156;
		#10; r229 = (8'h6d >=  ( ~ ( $time)));
		#10; r219 = ((r171 ? r116 : 25'h2ba2) | r103);
		#10; r178 = ( ( - ( (( ( - ( (r111 || r145))) ? ((( ( & ( r207)) + (r100 + (r85 / (29'h7a89 == 29'h73df)))) != (r191 === 30'h24b3)) >= (r163 == ((r136 % ( ( | ( (11'h78f &&  ( | ( (2'h1 >= ( ( - ( 10'h1d4)) > (7'h39 % 26'h14d3)))))))) + r43)) / ($stime >= r192)))) : (r211 === 10'h381)) !=  ( - ( 6'h1f))))) > (r63 !==  ( ~ ( (r71 / 15'h32a7)))));
		#10; r235 = ($stime === r52);
		#10; r181 =  ( ! ( (( ( & ( (r72 | ((r82 - (r122 - r110)) / 3'h1)))) > (1'h0 !=  ( & ( r117)))) % r35)));
		#10; r115 = 31'h222c;
		#10; r21 = 10'hbc;
		#10; r202 = (( ( & ( $time)) > ((r141 || (28'h91 ||  ( - ( 25'ha3e)))) || ((r78 & ((r252 >  ( ~ ( 2'h1))) > (r235 ^ $stime))) &&  ( & ( 9'hbc))))) == $time);
		#10; r255 =  ( & ( 30'h67f1));
		#10; r65 = 13'h342;
		#10; r208 =  ( & ( (9'h148 !== ((((r86 - r205) | 16'h10c7) + $stime) / (r145 /  ( ^ (  ( & ( 24'h4f19)))))))));
		#10; r25 = (r242 ? ( ( | ( (((((9'hab + (r120 & ((( ( + (  ( - ( r5)))) ? r90 : r232) % ( ( | ( (11'h6ec ? r150 : r41))) && 22'h5c1a)) !== ((12'hd86 * ((4'h5 + r76) * $stime)) != ((( ( | ( 28'h378b)) === 5'h11) != r235) >= 5'hb))))) != (((r232 !== ((r240 * r116) *  ( ^ ( (((18'h6629 < 31'h6fe7) * (28'h76b ^ 11'h18d)) > 32'h79d2))))) % (17'h4ad6 ? r19 : 29'h25f7)) | 28'h695e)) <= r176) !== 3'h2) === (9'h14f !== ((r71 %  ( - ( (r82 > ((6'h1b ^  ( & ( 22'h355c))) | 21'h4af7))))) !=  ( + ( (( ( & ( ( ( + ( $stime)) | r247))) <= 12'h5ff) | 5'h1a)))))))) < r124) :  ( + ( 25'h1324)));
		#10; r216 = 16'h6943;
		#10; r223 = $time;
		#10; r182 = r155;
		#10; r64 = (r73 - 31'h2134);
		#10; r254 = 9'hfb;
		#10; r180 = ( ( & ( ((r246 < (( ( ! ( r9)) <= r190) >= r25)) % (r150 != 6'hf)))) + 13'h1361);
		#10; r26 = (( ( | ( r12)) | r21) -  ( ~ ( ( ( ~ ( r129)) % (r99 < (r227 != (17'h1614 && ((r18 >= ((r85 % (r91 | r23)) <= 21'h2add)) === ( ( - ( r175)) === 15'h60cd)))))))));
		#10; r58 = (((26'h4eb6 >= r67) & ( ( - ( ((($stime <  ( ^ ( 24'h5968))) != ( ( & (  ( ^ ( r173)))) <= (($stime * (( ( + ( ((r216 > $stime) & r144))) || r153) &  ( | (  ( ^ ( $stime)))))) <= 22'h5feb))) % ( ( ^ ( r192)) +  ( + ( 9'h140)))))) | 16'h6670)) ===  ( ! (  ( - (  ( - ( ( ( | (  ( + (  ( + ( r128)))))) / ((( ( - ( (4'h3 !== r13))) | r212) >= (r48 + (18'h2621 != ( ( ! ( (6'h2b | r84))) / ((( ( ! (  ( - ( 1'h1)))) + r38) &&  ( ! ( r39))) == 21'h46a))))) != $stime)))))))));
		#10; r227 = 4'ha;
		#10; r151 = r208;
		#10; r180 = (((r193 || r112) & (r198 !== r202)) | r46);
		#10; r81 = (((r224 <= 27'h4c16) ? ((r96 == ((($time % (r59 && r245)) !== 28'h5b91) <  ( | (  ( ^ ( 22'h78)))))) + 30'h1c62) : (r225 < ((18'h2d37 < ( ( ~ (  ( ^ ( 25'h73f9)))) == 4'h5)) ? ((r158 & r216) - (r243 !== r243)) : 24'h2bb7))) > 1'h1);
		#10; r143 = r52;
		#10; r222 = (( ( ^ ( r10)) + (22'h3a15 && ( ( ^ ( r163)) < 4'h8))) !=  ( ! ( ((r119 % ((r184 || ((((((18'h62e0 ? ((r123 > r7) *  ( ^ ( r81))) :  ( + (  ( & ( r60))))) ===  ( ^ ( (2'h2 ? ((18'h261a - 14'h226f) !== (10'h88 / 25'h5b0e)) : ((16'h4605 * 22'h6ac6) == 14'h32ee))))) % ((r135 * 25'h303b) && 13'h143b)) % r94) &  ( ^ ( r16))) *  ( - ( ((((((r183 & r178) && ( ( ! ( 19'h2f4b)) * (31'h7e35 + 12'h73e))) > (((18'h5c0c === 28'hb1c) > (1'h1 || 5'h1a)) ^ r54)) ? r222 : 25'h54cf) | (r131 - (r248 & r78))) == 18'h5932))))) % r73)) < r194))));
		#10; r241 = $stime;
		#10; r4 = ( ( & ( r125)) <= (r41 ? ((23'h312d != r35) > r184) : ((19'h2838 + r31) == 25'h25bc)));
		#10; r65 = r4;
		#10; r68 = r86;
		#10; r46 = 2'h2;
		#10; r123 = ((((r247 || ($stime | r248)) ?  ( ~ ( ($time & (r73 === r43)))) : 5'h16) > 25'h4e87) == r2);
		#10; r177 = $time;
		#10; r15 =  ( ^ ( r236));
		#10; r236 = 25'hdf4;
		#10; r186 = ( ( ^ ( (r163 % ((r186 ^ ( ( ! ( $stime)) * $time)) && r104)))) | 21'h3b98);
		#10; r238 = (r170 + 1'h0);
		#10; r167 = r11;
		#10; r47 =  ( ~ ( (r164 !== (27'h2b93 | 19'h3f3))));
		#10; r152 = 13'h1ae6;
		#10; r136 = 11'h27f;
		#10; r87 = r50;
		#10; r44 = (r105 &&  ( ~ ( (((( ( | ( $stime)) /  ( - ( 21'h58a3))) * 18'h2973) > ( ( - ( $time)) ? (((15'h3f4c ^ (r180 - ((r233 * $stime) !== r28))) | 15'h4cb7) - (r234 * ( ( ^ ( 7'h4d)) > (((r200 && 23'h14a0) != r159) <= ((( ( & (  ( ~ ( $time)))) - r226) | 16'h45eb) - r22))))) : r232)) === r165))));
		#10; r85 = (r147 > r18);
		#10; r231 = ((8'h94 ^ 4'h5) ? (((r200 || ((($stime & r75) && 11'h0) & 32'h44a8)) || r49) -  ( ^ ( (r204 | r161)))) : ( ( + ( (14'h1ec9 ===  ( - (  ( & ( (16'h1ac3 == r40)))))))) <= (( ( - ( r196)) %  ( | ( ((30'h5eb9 | ( ( ^ (  ( ^ ( (((((15'ha3e + 3'h1) & r235) & (31'ha50 ^  ( + ( 21'h1246)))) != 4'ha) !=  ( ^ ( (6'h11 != r84)))))))) / ( ( ~ ( (r199 - ((((19'h6553 + 29'h2692) - 11'h87) & r215) != r247)))) & r129))) <= 10'h2d8)))) ^ (r63 == r161))));
		#10; r243 =  ( + (  ( ! (  ( ! ( ($stime >= r141)))))));
		#10; r225 = ((r227 ^  ( ^ ( (((r211 != r246) != 1'h0) / ((r151 / (r189 - ((2'h0 ?  ( | ( ((17'h15be != 25'h57cd) || r18))) : r130) <= r133))) > ( ( - ( r177)) & r100)))))) ^ (30'h29af ? r155 : r154));
		#10; r188 = r9;
		#10; r20 = 7'h30;
		#10; r47 = r47;
		#10; r58 = r172;
		#10; r25 = 14'h2732;
		#10; r120 = r209;
		#10; r234 = r122;
		#10; r109 = 32'h6179;
		#10; r220 = $stime;
		#10; r62 = 20'hf98;
		#10; r123 = 30'h434c;
		#10; r157 = ((9'hdf !== r221) != (r158 ^ 27'h7b5b));
		#10; r118 = r28;
		#10; r225 = $stime;
		#10; r144 = (r5 == ( ( & ( $time)) < ( ( + ( 19'h1ed0)) != 2'h1)));
		#10; r134 =  ( ^ ( 4'h6));
		#10; r6 =  ( - ( 21'h63eb));
		#10; r81 =  ( + ( ((((( ( + ( (($stime != (( ( - ( (30'h417 * 9'hd2))) !== (r98 && (31'h2b9b >=  ( - (  ( | ( 4'h2))))))) /  ( ! ( 21'h3fae)))) * r7))) !==  ( ! ( r89))) + (32'h6ea2 + r41)) % (6'h2b === ($stime - ((12'h589 || 3'h4) | (((31'h73e9 ? ( ( | ( ( ( - ( r222)) >= ($time + (13'h126a * 30'h491b))))) ? r80 :  ( ! ( ( ( + ( (20'h15ba >= 20'ha2))) >= (1'h0 === 32'h7b25))))) :  ( + ( ( ( + ( r171)) / 14'h2d54)))) === 20'h2b36) ^ r30))))) !== ( ( ^ ( (r242 - $time))) &&  ( | ( r56)))) * ( ( + (  ( ! ( 6'h35)))) >= (r1 - r197)))));
		#10; r156 = 18'h31e3;
		#10; r11 =  ( ~ ( r46));
		#10; r140 = r153;
		#10; r230 = $time;
		#10; r221 = ( ( ! ( 4'hb)) >= 11'h400);
		#10; r228 = 10'haa;
		#10; r125 = ((17'h2e5c >  ( ~ ( (r130 - r65)))) > ((r27 - (((r7 ==  ( | ( (((r242 ||  ( ~ ( r127))) *  ( + ( ((((r163 >= (18'h76bb == 3'h1)) & r140) ? (r137 == ((19'h1a8 && 20'h4b97) == 22'h44f5)) : r210) ? ($time / 23'h2b69) : r56)))) <= (16'h5540 +  ( ! ( r90))))))) !== r76) &  ( ! ( (r21 < 31'hbd9))))) + r248));
		#10; r160 = ((25'h1e99 &  ( - ( (((r104 & (r27 | (((17'h320e || r91) - (r111 != 31'h23ab)) !== r116))) % (( ( ! ( r132)) <= 21'h7a3d) || (((r78 != ( ( ! (  ( ~ (  ( ! ( ( ( ^ ( 8'h8)) != 3'h6))))))) < ((((r197 == $time) +  ( | (  ( ^ ( 17'h4d54))))) && 6'h9) -  ( ^ ( (( ( ! ( 7'h48)) %  ( ! ( 8'h7e))) != (24'h38e3 || r47))))))) + r108) >= r183))) ^ r103)))) && 20'h1ff0);
		$displayb("r0 = ",r0);
		$displayb("r1 = ",r1);
		$displayb("r2 = ",r2);
		$displayb("r3 = ",r3);
		$displayb("r4 = ",r4);
		$displayb("r5 = ",r5);
		$displayb("r6 = ",r6);
		$displayb("r7 = ",r7);
		$displayb("r8 = ",r8);
		$displayb("r9 = ",r9);
		$displayb("r10 = ",r10);
		$displayb("r11 = ",r11);
		$displayb("r12 = ",r12);
		$displayb("r13 = ",r13);
		$displayb("r14 = ",r14);
		$displayb("r15 = ",r15);
		$displayb("r16 = ",r16);
		$displayb("r17 = ",r17);
		$displayb("r18 = ",r18);
		$displayb("r19 = ",r19);
		$displayb("r20 = ",r20);
		$displayb("r21 = ",r21);
		$displayb("r22 = ",r22);
		$displayb("r23 = ",r23);
		$displayb("r24 = ",r24);
		$displayb("r25 = ",r25);
		$displayb("r26 = ",r26);
		$displayb("r27 = ",r27);
		$displayb("r28 = ",r28);
		$displayb("r29 = ",r29);
		$displayb("r30 = ",r30);
		$displayb("r31 = ",r31);
		$displayb("r32 = ",r32);
		$displayb("r33 = ",r33);
		$displayb("r34 = ",r34);
		$displayb("r35 = ",r35);
		$displayb("r36 = ",r36);
		$displayb("r37 = ",r37);
		$displayb("r38 = ",r38);
		$displayb("r39 = ",r39);
		$displayb("r40 = ",r40);
		$displayb("r41 = ",r41);
		$displayb("r42 = ",r42);
		$displayb("r43 = ",r43);
		$displayb("r44 = ",r44);
		$displayb("r45 = ",r45);
		$displayb("r46 = ",r46);
		$displayb("r47 = ",r47);
		$displayb("r48 = ",r48);
		$displayb("r49 = ",r49);
		$displayb("r50 = ",r50);
		$displayb("r51 = ",r51);
		$displayb("r52 = ",r52);
		$displayb("r53 = ",r53);
		$displayb("r54 = ",r54);
		$displayb("r55 = ",r55);
		$displayb("r56 = ",r56);
		$displayb("r57 = ",r57);
		$displayb("r58 = ",r58);
		$displayb("r59 = ",r59);
		$displayb("r60 = ",r60);
		$displayb("r61 = ",r61);
		$displayb("r62 = ",r62);
		$displayb("r63 = ",r63);
		$displayb("r64 = ",r64);
		$displayb("r65 = ",r65);
		$displayb("r66 = ",r66);
		$displayb("r67 = ",r67);
		$displayb("r68 = ",r68);
		$displayb("r69 = ",r69);
		$displayb("r70 = ",r70);
		$displayb("r71 = ",r71);
		$displayb("r72 = ",r72);
		$displayb("r73 = ",r73);
		$displayb("r74 = ",r74);
		$displayb("r75 = ",r75);
		$displayb("r76 = ",r76);
		$displayb("r77 = ",r77);
		$displayb("r78 = ",r78);
		$displayb("r79 = ",r79);
		$displayb("r80 = ",r80);
		$displayb("r81 = ",r81);
		$displayb("r82 = ",r82);
		$displayb("r83 = ",r83);
		$displayb("r84 = ",r84);
		$displayb("r85 = ",r85);
		$displayb("r86 = ",r86);
		$displayb("r87 = ",r87);
		$displayb("r88 = ",r88);
		$displayb("r89 = ",r89);
		$displayb("r90 = ",r90);
		$displayb("r91 = ",r91);
		$displayb("r92 = ",r92);
		$displayb("r93 = ",r93);
		$displayb("r94 = ",r94);
		$displayb("r95 = ",r95);
		$displayb("r96 = ",r96);
		$displayb("r97 = ",r97);
		$displayb("r98 = ",r98);
		$displayb("r99 = ",r99);
		$displayb("r100 = ",r100);
		$displayb("r101 = ",r101);
		$displayb("r102 = ",r102);
		$displayb("r103 = ",r103);
		$displayb("r104 = ",r104);
		$displayb("r105 = ",r105);
		$displayb("r106 = ",r106);
		$displayb("r107 = ",r107);
		$displayb("r108 = ",r108);
		$displayb("r109 = ",r109);
		$displayb("r110 = ",r110);
		$displayb("r111 = ",r111);
		$displayb("r112 = ",r112);
		$displayb("r113 = ",r113);
		$displayb("r114 = ",r114);
		$displayb("r115 = ",r115);
		$displayb("r116 = ",r116);
		$displayb("r117 = ",r117);
		$displayb("r118 = ",r118);
		$displayb("r119 = ",r119);
		$displayb("r120 = ",r120);
		$displayb("r121 = ",r121);
		$displayb("r122 = ",r122);
		$displayb("r123 = ",r123);
		$displayb("r124 = ",r124);
		$displayb("r125 = ",r125);
		$displayb("r126 = ",r126);
		$displayb("r127 = ",r127);
		$displayb("r128 = ",r128);
		$displayb("r129 = ",r129);
		$displayb("r130 = ",r130);
		$displayb("r131 = ",r131);
		$displayb("r132 = ",r132);
		$displayb("r133 = ",r133);
		$displayb("r134 = ",r134);
		$displayb("r135 = ",r135);
		$displayb("r136 = ",r136);
		$displayb("r137 = ",r137);
		$displayb("r138 = ",r138);
		$displayb("r139 = ",r139);
		$displayb("r140 = ",r140);
		$displayb("r141 = ",r141);
		$displayb("r142 = ",r142);
		$displayb("r143 = ",r143);
		$displayb("r144 = ",r144);
		$displayb("r145 = ",r145);
		$displayb("r146 = ",r146);
		$displayb("r147 = ",r147);
		$displayb("r148 = ",r148);
		$displayb("r149 = ",r149);
		$displayb("r150 = ",r150);
		$displayb("r151 = ",r151);
		$displayb("r152 = ",r152);
		$displayb("r153 = ",r153);
		$displayb("r154 = ",r154);
		$displayb("r155 = ",r155);
		$displayb("r156 = ",r156);
		$displayb("r157 = ",r157);
		$displayb("r158 = ",r158);
		$displayb("r159 = ",r159);
		$displayb("r160 = ",r160);
		$displayb("r161 = ",r161);
		$displayb("r162 = ",r162);
		$displayb("r163 = ",r163);
		$displayb("r164 = ",r164);
		$displayb("r165 = ",r165);
		$displayb("r166 = ",r166);
		$displayb("r167 = ",r167);
		$displayb("r168 = ",r168);
		$displayb("r169 = ",r169);
		$displayb("r170 = ",r170);
		$displayb("r171 = ",r171);
		$displayb("r172 = ",r172);
		$displayb("r173 = ",r173);
		$displayb("r174 = ",r174);
		$displayb("r175 = ",r175);
		$displayb("r176 = ",r176);
		$displayb("r177 = ",r177);
		$displayb("r178 = ",r178);
		$displayb("r179 = ",r179);
		$displayb("r180 = ",r180);
		$displayb("r181 = ",r181);
		$displayb("r182 = ",r182);
		$displayb("r183 = ",r183);
		$displayb("r184 = ",r184);
		$displayb("r185 = ",r185);
		$displayb("r186 = ",r186);
		$displayb("r187 = ",r187);
		$displayb("r188 = ",r188);
		$displayb("r189 = ",r189);
		$displayb("r190 = ",r190);
		$displayb("r191 = ",r191);
		$displayb("r192 = ",r192);
		$displayb("r193 = ",r193);
		$displayb("r194 = ",r194);
		$displayb("r195 = ",r195);
		$displayb("r196 = ",r196);
		$displayb("r197 = ",r197);
		$displayb("r198 = ",r198);
		$displayb("r199 = ",r199);
		$displayb("r200 = ",r200);
		$displayb("r201 = ",r201);
		$displayb("r202 = ",r202);
		$displayb("r203 = ",r203);
		$displayb("r204 = ",r204);
		$displayb("r205 = ",r205);
		$displayb("r206 = ",r206);
		$displayb("r207 = ",r207);
		$displayb("r208 = ",r208);
		$displayb("r209 = ",r209);
		$displayb("r210 = ",r210);
		$displayb("r211 = ",r211);
		$displayb("r212 = ",r212);
		$displayb("r213 = ",r213);
		$displayb("r214 = ",r214);
		$displayb("r215 = ",r215);
		$displayb("r216 = ",r216);
		$displayb("r217 = ",r217);
		$displayb("r218 = ",r218);
		$displayb("r219 = ",r219);
		$displayb("r220 = ",r220);
		$displayb("r221 = ",r221);
		$displayb("r222 = ",r222);
		$displayb("r223 = ",r223);
		$displayb("r224 = ",r224);
		$displayb("r225 = ",r225);
		$displayb("r226 = ",r226);
		$displayb("r227 = ",r227);
		$displayb("r228 = ",r228);
		$displayb("r229 = ",r229);
		$displayb("r230 = ",r230);
		$displayb("r231 = ",r231);
		$displayb("r232 = ",r232);
		$displayb("r233 = ",r233);
		$displayb("r234 = ",r234);
		$displayb("r235 = ",r235);
		$displayb("r236 = ",r236);
		$displayb("r237 = ",r237);
		$displayb("r238 = ",r238);
		$displayb("r239 = ",r239);
		$displayb("r240 = ",r240);
		$displayb("r241 = ",r241);
		$displayb("r242 = ",r242);
		$displayb("r243 = ",r243);
		$displayb("r244 = ",r244);
		$displayb("r245 = ",r245);
		$displayb("r246 = ",r246);
		$displayb("r247 = ",r247);
		$displayb("r248 = ",r248);
		$displayb("r249 = ",r249);
		$displayb("r250 = ",r250);
		$displayb("r251 = ",r251);
		$displayb("r252 = ",r252);
		$displayb("r253 = ",r253);
		$displayb("r254 = ",r254);
		$finish(0);
	end
endmodule
