/*
 * Copyright (c) 2000 Stephen Williams (steve@icarus.com)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 */

/*
 * This test checks that times within modules are scaled up to the
 * precision of the simulation.
 */

`timescale 100us / 1us
module slow (out);
   output out;
   reg	  out;

   initial begin
      #0 out = 0;
      #1 out = 1;
   end

endmodule // slow


`timescale 10us / 1us
module fast (out);
   output out;
   reg	  out;

   initial begin
      #0 out = 0;
      #1 out = 1;
   end

endmodule // fast

`timescale 1us / 1us
module main;

   wire slow, fast;

   slow m1 (slow);
   fast m2 (fast);

   initial begin
      #5
	if (slow !== 1'b0) begin
	   $display("FAILED");
	   $finish;
	end

        if (fast !== 1'b0) begin
	   $display("FAILED");
	   $finish;
	end

      #10
	if (slow !== 1'b0) begin
	   $display("FAILED");
	   $finish;
	end

        if (fast !== 1'b1) begin
	   $display("FAILED");
	   $finish;
	end

      #80
	if (slow !== 1'b0) begin
	   $display("FAILED");
	   $finish;
	end

        if (fast !== 1'b1) begin
	   $display("FAILED");
	   $finish;
	end

      #10
	if (slow !== 1'b1) begin
	   $display("FAILED");
	   $finish;
	end

        if (fast !== 1'b1) begin
	   $display("FAILED");
	   $finish;
	end

      $display("PASSED");

   end // initial begin
endmodule // main
