module test();

reg [0] illegal;

endmodule
