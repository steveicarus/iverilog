module test();

parameter name = 1;

endmodule
