module module_0 #(
    parameter id_1  = 32'd92,
    parameter id_3  = 32'd50,
    parameter id_4  = 32'd25,
    parameter id_8  = 32'd99,
    parameter id_9  = 32'd40
) ();

  // Cannot assign to a parameter.
  assign id_8 = 1;

endmodule
