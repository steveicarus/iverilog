module test();

reg [] illegal;

endmodule
