// Check that declarations for dynamic arrays of dynamic arrays are supported.

module test;

  // Dynamic array of dynamic arrays
  int q[][];

endmodule
