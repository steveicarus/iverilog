module test();

typedef enum { a, b, c } enum_type;

enum_type enum_value;

initial begin
  enum_value = 1;
end

endmodule
