module test;

wire [7:0] value, value;

endmodule
