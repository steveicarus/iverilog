-- Copyright (c) 2015 CERN
-- Maciej Suminski <maciej.suminski@cern.ch>
--
-- This source code is free software; you can redistribute it
-- and/or modify it in source code form under the terms of the GNU
-- General Public License as published by the Free Software
-- Foundation; either version 2 of the License, or (at your option)
-- any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program; if not, write to the Free Software
-- Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package vhdl_range_pkg is
    subtype integer_asc is integer range 0 to 7;
    subtype integer_desc is integer range 8 downto 1;
end vhdl_range_pkg;

package body vhdl_range_pkg is
end vhdl_range_pkg;
