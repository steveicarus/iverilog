module test();

parameter y = 1;
parameter a = 0;

parameter x = y ? a : b;

endmodule
