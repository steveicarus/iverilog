module d();
       nand n2(w1,

       nand n1(w2);
endmodule
