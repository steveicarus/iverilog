/*
 * Copyright (c) 1999 Stephen Williams (steve@icarus.com)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 */

primitive BUFG ( O, I );
   output O;
   input I;
   table
      0 : 0 ;
      1 : 1 ;
   endtable
endprimitive

module main;
   wire out;
   reg in;

   BUFG #5 bg(out, in);

   initial begin
      in = 0;
      #10 if (out !== 0) begin
	 $display("FAILED -- %b != 0", out);
	 $finish;
      end
      in = 1;
      #4 if (out !== 0) begin
	 $display("FAILED -- %b != 0", out);
	 $finish;
      end
      #2 if (out !== 1) begin
	 $display("FAILED -- %b != 1", out);
	 $finish;
      end
      $display("PASSED");
   end
endmodule
