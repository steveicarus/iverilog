module top;
  buf(strong0, highz1) #1 sclbuf0(iscl);
endmodule
