// Check that an error is reported when trying to bind an argument by name that
// is also provided as a positional argument.

module test;

  function f(integer a, integer b);
    $display("FAILED");
  endfunction

  initial begin
    integer x;
    x = f(1, .a(2)); // This should fail. `a` is provided both as a positional
                     // and named argument.
  end

endmodule
