module test;

// synthesis translate_on
// synthesis translate_off

initial $finish(1);

endmodule
