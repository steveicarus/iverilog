`timescale 1ns/1ps

module top;

  initial begin
    $sdf_annotate("ivltests/sdf_header.sdf", top);
  end

endmodule

