module test;
    initial begin
	$mytest(1,9.6,3);
    end
endmodule
