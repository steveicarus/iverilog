module test();

typedef enum { a, b, c } enum_type;

enum_type enum_value;

assign enum_value = 1;

endmodule
