// Check a missing local time precision.
`resetall
module no_ltp;
  timeunit 1ns;
endmodule

