// Check that declarations for queues of unpacked arrays are supported.

module test;

  // Queue of unpacked arrays
  int q[10][$];

endmodule
