initial #1 $display("PASSED");
